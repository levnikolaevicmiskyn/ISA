caran@LAPTOP-FP3DTT1V.10520:1608453886