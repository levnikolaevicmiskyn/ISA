../../../auxilliary/dadda/MBE_24bit.vhd