../../../auxilliary/dadda/MBE_32bit.vhd