GIF87a��     ����    ��� � ����� KKK���������������������,    � ��I��8�ͻ�`(�di�h��l�p,�tm�x��|����pH,�Ȥr�l:�ШtJ�Z�جv��z��xL.���z�n���|N�����~������������������������������������������������������������������������������������������������������������������������������������ 
H����*\Ȱ�Ç#J�H��ŋ3j�ȱ�Ǐ� C�I��ɓ(S�\ɲ�˗0cʜI��͛8s��ɳ�ϟ@�
J��ѣH�*]ʴ�ӧP�J�J��իX�j�ʵ�ׯ`ÊK��ٳhӪ]˶�۷p�ʝK��ݻx���˷�߿�L���È+^̸��ǐ#K�L���˘3k�̹��ϠC�M���ӨS�^ͺ��װc˞M���۸s��ͻ�����N����ȓ+_μ���УK�N����سk�ν����ËO�����ӫ�����(���>{��'ط�?���������I0��' �	�g��&���:��68�Z�!�nء�f(!�(b�+��b�*�hb��`��b�5�x��#�xb�3�H�C�h�~BҨ��Lɢ�.$�<>Yd��Y�ޗx)��`�y�ud��e�j��n���r�y�v��hx���n}�)�m�jhl�:]��6���FJ��V���f��Z�n��d�~*�c��jjb��
(����j�ϥ�����j�sފ�r��&� �+�`��&����6���F+��Vk��f���v����+��k�覫��[-���B���*��Pl�L0�� K��0���p��0�/q�W,��_�q�O�1�or� �,��$��r�,��2�/�s�0�,��4߬s�<��3�?�t�@-��D�t����� �ދ���Я��o�K�5�_w��b����a�M��f����o���r����q�M��v�7�\o���'P�ۯP|u�����~C.���my���c~��gι�.��wnz�/����Ϋk	�&�/֋�>������~���.|���>����<��^�5��[�+�SOx��+�}��c����>�ݓ/~�㧏>��R�8Ԅ�`xn�ʋ���k���������[_� H@p�, �8��.j�+�������i̠5��.��ܠ=��0��s�����)v�	MH�ڰ�8D�i���0�<�\���MPj������C&��P|�HE'V1�W�\��*���I�MC��Xh�2bьSDcר�6��iT^ǈ�ƯL���V�A8�яn�� �8�@�L����/JMMy����WH@Z���D�%5�IEvr�4����Y�}��$'W��V�򕟌%+a9KJ�r��L��w�^�ҕ��%0g�b���_{�?J~�񂗻�I�jZ��̦6���nz���8�Mx��L^$�:��+���u�d��8�u���K����F��L@�O�����$�z�gρ*��oi�=��{!t��([*�\Z��̨Fղ�x�S��1eG�9ҸԤ���HPҁ��-5�J���7�i�z�ӱp��)mzϢ�����t)T�:�-/�)Q3���0�u��[vP�JO�d��XIZՆ�U�Tm+Kך��Jt�読>
U�j����`K�����M�b��i���*F�ꪏ��Ѥ]M�)��3����gC��m�yz�@Z�J��&�}e-v)8f�����-iw;���ַ,[f3��Y�ε�3�j1�{�S:.����o�]�J��T\�s�;���3�]��j9����轮z��^�׽%�&�ڴ�5L�nX��>�.��mo��K��.��v+Y����u�d�Y\��VFp�7\`w��^�py����oE���{��2N^�q�e��۸�~Ta#��Z�z1� 5�l[<���� �q��Lc&#�����-0�z�v�(f��4�6��O���<f1k1���r��{_����[���Gf'���v�s����Q�n��㯏�l����z/~.���h33Zώ�t�tlG�6��������I�Ѡ�t�MjI��b��qd�KY�d٤qF�f�l�R��ָ����yZ�v��ms"ܜ*'��t wm�S7�ٹvv2��E:�y�@��W�X�5������M�r��܄�vM�ca�'��^���MW��تeu����
��/yuT��Rzk�� �0��cה��d\�}i���61�o�X�r�8�'ro�f��S�e�����#_��O�c6�:Vh�w�����\�fx�J�[��)�8�9.�Ey\�&�7�MRr�F]��u�e�Np��|���Mk^�lW�R�8�����<�f��Ra^�~���/.��s����X��H��b*����ؿ+��#��/��ܳZ��'������F��Ι��{���wD�m��C�t�^=�o��Aۋ�|9��q�m{����Ϻ�;�����#n�6�OO����G~�I���k����}����|�L-�+�����~������-�bA�X�����������Ͽ���mz[� �/�n_gyhg?h�Y�`��G��l�m8��>ƒ4�_L����H�'^$�K(3bFV;^3"(��*��,؂.��0�28�4X�6x�8��:��<؃>��@(�seE�KC��e{G�~�N��-�TX�Vx�X��Zh-S�-�`?�n�w�'h�q{����>�rx&��� n `8pH'db�\%�oh у�s(Ay�T�hD��WsȆ���H��F��H��x&~���(��Ј�B �0�h�}���*o��]��Z�A��x��H������!������2�������%
��ȋ������H!�� 2⋰��Ѹ����ڨ��H���������⍸��x����{������Q�꘎� �x�و$�������8� I����H��ȉ�Xh�Ww.W��Ax)Gg(?���R �x�+�%�H�ző�5�x�����_䋅c�o��S�����y���6��ؒ6I��8���@����}'G|�~Z��~Be{�H�����x5I��8���������8��莯�<9�凞���X)�Mɕ��/kY�b�0��f�3����i�d��Ԉ��ؗuI�lY��蕃�������i��y��P9{�u�gS��T�,�@���;i}f���y�bx�Y�Ip��ؘ�����Q}����|�p���\FYY�pEt�tշ��)�T��������ȍ�Șx��wi��h��	��I��G����o��I�{���ٔ�)��X���	��	��I�ڹ�����	��y�C�T�z�w�W��Xy�)y�y�b�})[���10���S����ڡ����:�$Z�&z�(J�J�49[��Qg�{y�+J�ɠ/ɢ*&�i=
�@�R�	:?�(T����|2������r��w����R ����Y�빞[Y�$I�����y�[��p�P�O�yy!*`z�z� qJ�{��
 zJ��ʧ�X Wꆅ�q�{�]:��5RJ�
�cz�� �`�`��W*�툝�R��sz�����ʖ�Z�4E��w��u�H�h8�"p����FڛΘ����zA"�:Z�d�U�h��y�)�����!*�n�ؚ�ڊ��j��J�������)�źc��/�ح+���薂����S@g�
:tX���א����^ԗ���o��
��۰�: {&b؟vH�+{!��-����-�9��:��*�s8-:9��ʧ
.��?��;������
ɤ���j�x!0��U�������z���J��k,
+��myG
k!Ω-�W�-�)��*0�B�������H�i��A�z;�}p֚���ɹ{��2��V*�5���Z��*�|D��
��X�����B8��4�ʷ��4�����<�۩�*��K��+�ĩ�Z�s���J��K��:�{��ظ�{A�#�����:��K�#۷�˗����
�?+��G��j���J��zEۚ�+�7zSQk�B	�����ڑi������������y�IU�PK����L��K�4I'���
��k+��;��W��W�Se�釜��L�h rh ����l��� |�;�K��X���S������+ L��Vy��X���X�䩻�[GMi����j����8�D\����8����
�vX��� &�)l�+ Q,�,+l����;&|&[L�Yl�-��]����2l�KI}	z�!��J��j�e����}�ǂ\�&L�g"��۶�j�љ��[e,A��!i��l'��X������7���!������&�FȁL�\Ř+�5ڢ�-�	Yl��8Ő,�d�˾�˽̃�C@'��Ǭ��¬�����ǀ��|v
ɳԫ���SL�V��sx�Z��f�2Ť;ƦK���/"�΂���j��Β\S���I�����P <����i��КK���,��*��z�e:±{� ܩU�����/eܺ����3���M��|����q|���̓���-�j<�2]�ͻ���0��,���A��7����Ȋg�v���[����
�=���˫�@]Ɇ��w���ȵ���|S�<;�<�Hm����&���m����ۢK{�D5U}y��x�֣���R�ؽ^}����X-̫\�V�ˈ]��׼|Ռ��3��O����,w���g�m��;}�Y��U\���)��#��ֹ�",����,-L��Ħ
�1\��Vb��S�JL��zõm�BL����A��(L�;M�0�n��o캾�����D�7+ï�<�3��h����ѓ�ݻ�����f�ŧ������o<����y��>�ا�����l��L��ڽ��vL�I*֑M��<����k�q��S���gxn�0�i-�,���� ٴ��;�����6�Gk��ZՒ����k��W������-����Z���P=��q~]7ǌ��?]ݬ=�W����{;ߴ�ΉY���ݿH���B}�L<���/\�=���	ͥ�XS=�Ѣ[Ѻ�Ӈ�ї=�Q;�~��.|�ٸ�����m�ln��Cm݂�?���������B��EM�G��>�g��$���S��Y�������K�ȣ��LSw��V<̮̂�c������;��)��"��$>׻���~����F�����5މ�n����������ƴ��C��0���.�K�뙝po'Չ�b��u�|]��[lږ.����؝��m������������Z�����h^�ம���]�ɸ�r=����b�g��_^��>��Ѝ�o-����3^޼l����[�՛��ם�n��b����9����B��>o���J�TzW��{}�޾�\���칎�+�����޾(^��>�*����͎�.Z�_O^�e�Kz���3��ߺ�������a��D��x<�n�xD��Ι�&��t�����2F �n��Մ�Ȣ��oMN��G�"��_����M����ׅ�ҙQ?Q������lF�3�1 ���������S(��?���Ɵ��Z��O�Ώ���ϟ��O�(=�՟��?F������k��/����%�?���?�џ���տ����?��UN����ϩ����o�0�b�;ޚ/�ƮɳCE�M�5vٴ�o���y�{�.�� ���D*�K'�$�J���v����{�gtZ�f��ox\>���w|^����ƻ0A�16-�-+ī�ƨ&H @�H�J'@Kʍ#�&#��GJRKN�QM�T�ʬ,��(�����\�]�^]��UZ��K0QQYTc���楀)��d�W��UIG�a����hf��Cr�G�S�аp���%��J���s�b}�g���'�`A���)��/X�R�$"*��ʠ���l����G�!E�$Yr�:[0�a�&��,dΤY�&�7u���ӧ	�A�%Z3[Ѣ��.��ԩL-V�<���թ7ab���W�1��K6�X�W�VU���[�q����u��6�V^ă��_��&\���1{ɔI���9F&MVB�S�N�%U��Y�Ϙ/g��t�ӢM�-��Μa�1rj�ǶLH�[3�^�{��;Sۚ��Ǽ�NԼ�O�$��ە�o�>�z�s⬳S�lz�q��7{V�}�i��ɯ^�������?_v<��h���%:�BlAt�A#ı/ ;C%Y�0����T����
s���
|/�,DL#�#p����H3>�C�.NL'�w8�q�'��Q��,Q	\(�/��ыԛ2 �$D#�q�.��ѥ�`tC���04Ѵ�B-:Pþִ�N<��s�<��%:3���3�������
�Ͽ�\CF�`qT)���L�pL�R��sm�c u�,�.��QV�9�P�F�tV_F;�?�@��;SaM:�`H�O�ݴUcMMYe��M@��А@5�L>��v[n�=l�j��2\�ԣM�Ԉ�%�3D3��֋8����r��W{}��]6\U�$��[6���Z#��.0��5]~��ې�D���pq96�d�SFy_|�,�����5��v�Y����{N�f-حggS�wٙWU����+:��+�X��:�X�6^�g��n�.�,�<��Mi��v�Y�ac9^�G��|�U�{o���pnz�|\
I<Wc��M����7p��h��1Y��Z�+_c�q7ޜˋ|3��G�k�w��[�s��1\PZ��p9�34�6S�i���S\t?7�x��(sG6p�g߱��L��V��������j�?�m�:4_5k��gs�>J'I�{��7��
���~MYu��h�V�(�g~����ާ�P�ܣ�� �� 9/f�r��<�A��uv �G����N�KS���1�u�q[Tʐ��)7�S��f�R�.x�cC�$fC�e�u�]�r'L����dl��2Mu-d��A	f�#!��9�P�kdc����f)�]��v��}��ѨcD_��<��ȧ=<�&�{d��v���*}�)׼W����� d$���8-{�A  y��F��z�`*-XAA�cq��舆�Q����H8��χ�ca�(�\�� В�p�N�b_8����C/���Y� �E"n��]���Y#*Yi���ar��*)�\V\�9�����!K�.����r��f-���^&T��C2�=Z�2i<}��F�5�4%/�c��X�|X;���Үŧ��z��N��d+�V���ÒE�Z/4K��N��S�����J�EP�S�i8%gBp*��chW��U�"Ɍ�+(B��8.hU]�RX�Ğ*�_K��"�9��"�6,��J��pr_�O���vb�&A�RF%�FV���le�I�3��b�^^��U��V�^uh��gK���kgS�Z\��*�V��nUT��8ȡ��j�:f�e�ג�9��J�����*|=�OT�c��$G�0p�svB+fZV����ԗR�7�P��,�z�9�q��e���'v���+&�8O�@�]0 �˅������_��U�  �J`P���EՄ�5�� Fw��k�!4�Q<X���D��F��K�5Q�0�&GE��s4f�	@�����ð�n����Y��&E�������1��f����WHq���e��/p�l���mv�X�l��;���Y�,-j9x^5N��%-��P�[�������g^������۳�mj7��X-M$k`�]�2�SK����_@�x3�5�e#hB�-���"�а����0t˴�C76���4$j)�˓��+lSw�v��C-մQ��v��V�:glg{ou>hc�;=��И���R=�)Z��0^	T�$	������IN�|��V�B��fۗ�ت{��]�Ȇ{�Ø|k�nH%'��-{���w�;�b�����]�@�:Vϲ��o�v�]���Z_�&�Wk=���>��)�����Tt��vH�V��GkrP�}�z�h���35I�`2�����@E喩�h���<F��kg;pr��+S�5�1�l��F�]�{M�wI�دl���ӊ.�~y������xlf|�o�i,��J"���I�@Kv��r�eǩ�KD')�(L��[�7���A�cs�
�z��
u>8��+��@�����sRI5Z"��/�L�9���D'f.k�*� 3z��yNC�H~�VcK��}�$Ͳ����/w^�cn��]�f�09ד�`�<8{<L@��ū6<�0=�̫��/F	4�5��+S�EK��(:�ɔ(3<�(���G��-����4��´ܨ���4T��X�@Q+��S6>��� �	j4���[B&��@_�A����(6���c�eS6�{��5��Ԫ<@<C4n3@�I#mJ�û�<5��"ᎏ�R�0��B`= �!���/����C�=���!��@#�BS�J�2��7%$۫��Ҁc*Eґ%B;��s�|9��A2��EZ$���8�;@��i����oJCa�;���@/�X9���[���#�"�;R���P�\�&,0� Ef�Ad��;�0:M�Ơ��rD�+P��5�[��YG�:5�@� 5�����邸�1��9*P�$�h�"�Q,.x�뮀�3#|;�x�L)���;$6�ػ3�H/B)�B�s���2��1-b|�I�d�p�����������ڃ�<��0��/�+0���4�{��K7�QĒ��;�Ct�v���I*��:j7n�7����?z�5��?�ѣ>�#��<.r���僺�<.R����-G����3���Lȝ*B�(�]�64�X�20�?�C0���C������F�z3��I�Ϳ����������
��.�p��0��$�&�͈�+��M�l��0�ߜ,ܔ���M�\��h��4
�	Ɋ��M�|M�Ν�pM��
�\���	�TF$#M�,O��0H�|5��
d�WK����8cx�O����|υP��9Y���Z�����\P�cZȼF`�s3��8	��D��
Uc�m`��$xFG�P�PH�8q��|���O5 �/�������e� M�����8�4O$M�l��kR�`����Rx�Q��0HQ"����	 �,eX8-p4���3űA�R0}y���0� 8-S=���������<��]X:u1T+��5�S� T��Sh�2�����PM�T_�	I�T=��`�Vp)��(��)U�#URW}��2M����
��
����|��B�����`�	au�҃�����MՔ��<�ӬMZ���Uk��]M��<N^u��V��b5��tN���f�UT�dmW� q�딑b�w��K= �|y�_�U-V�?�(���שج��v�b}�'V�����=X����Xb��a]M��Ul%�\�[�N��U�|�U�mYB� �k��;+Jۙ�0��-tt�[!�Hi�ۈ�s��B��:�x��$�����0)���Z���G:�1%�t:m,�Q�#l:Hu��E�dYG)��|][N}�M-Z��3�k8�<�ZI��[��!8(�9iCri���I���_dHm����E���Q\�%ސ����(������)&����\/L,��u�V֬	\� C�D�ͽ�ˡ�� ��5�j�ܓ\�C��G���SݐJL�D}q�=����I�M�54#��U��̾�^$5F�Q�d�oTA�U$�24 ꚜ]���\�=��%/�g��C ��ӣ��N���������	�iZ�}�`�8���%�� �]옺[`�])
��[��Z��F��W ;���/�i��=1g�#�����6�a%���I6L8����pl(�u�.��֥Cک�x���_!�(3����k܆rZ)�)>]�u��s��Zo�ax+L�\�8�!7�\ܹ����\������ �&���RdނY^��p^(�����$@��a�aE&χR���:е��B�[��w��Cx���ż2��`��\�����d+h0v��B�m�!1�}eY��B)��ɲi�G#�W.��mF�`�(�bޮX��a�䈻>���P��I7�;veH���zH��^�[i��^dr�3����I�����7ֱ�!�� .��&=�c9��e9υB�{	[R��1�"���b�k3";��$�|��F,c�8�0��@�|=�](f�����ʥ=f�A 1�}�᭡l}Թ^r7� d�Fz����2�r�i�T�p��gΨ{̤�u��B_�ڞ|lBr5���_۠�����c�`�:S֚���G�|˹��¨E��(F���ȺTc� }Eݡ됾ЮeZ�h��`z���=I�*_F����ij9�^���a�<7<d�Nd��e��1����l*�e��M�؂����ɢ��&h@�hƓ��m\���@�.v�+��Ж�����=�V^sC�c�k���.Y���ԃ����m#d�:�q��yM���7Фl�F@������\i��]�+�V� ;� �e�Ò��&�Q���	���oo�&�䞺��܍���� �KLy�d����D��5��)��E:���y|��*I+)Q�衕��>���َ6��#q����f��b��o�m�^G�p�kF��f�
���f�v���r��Y��aC���Tc�ė��B�=Q�+y*���m4�T��5ņA��M��+�H��/v5��E\޻�/�=MĆ�k��qwvk��p�5c:ǹ�K�F�/s�k��Rh��i3��魛t��u�rT!���Ȗr��%��P�-�0'*v�s\f�N�N����|<����
t����ZN-�
� �>�,[�0W?�B�Dq�Sj��K��St%���ptHOr��s\#�&��I�7���}lG��$�j�U?F���Nu�!���&u�d�)���K"{����ⴲs�=^��ʸ��I�ry�C+����]@�����)'�p�eBj�2f�h@���!t�T��EtCw����킚�s%[0�q���-�!�-�l���r!j(���-����쀯�߉�r~�@��]`��dq�[F��J0;!��|��`p���!d'�fb����Ӓ+�{i0fp�&������ѝ�,�娒8���k��>Nz'
�cP�g��ѕ��y#������?q��K���q���ݸ��?�D)��������zO;1do<f�P�z��Q/����S�g8����%�o3cmV��x�x�k��"�{�b]&y�g���5���:�t�a�/1��=����P�?�q?L��8L ��}m�]B��$��+�y!	�[k�X�ߍ�!�	.Ґ(�,g�g��I��R���f��-�k����3:�^���7<.����{���|q[�S��������⌈�ˊL�#c"#_@LK�!_A��(i��)*�d��@cd�&G����f%��-c�A�pj��1r���m�%+N��Ha�'ɮ� �@n�/����I���@FŁ�G{{KN3#�I�@>���o�!:u���r,����#?z�|0��GED� `��䣧~e�X�0�8 �!�OK5z�Ьi�&Μ:w���s��y/]Y9P6�\&��M�MDo�H��*2I[Ii����Le�U��@0	Xײm��L�^���
�a ,]�ވ��I��I� �%��@������4Ԉr��E�s�a�#Л9�p�#��"Q�<��B�Ѩ�i�6�ܺw���4Nk�e���}&��[����jy�D���̂��#�-W����~�9bJ{���8�K>�kB���j����ay�Mr�t���8��d�F�pB�]�Q2�?&�Ê<�}7�.PA6R V��=�������,�ނ��\���I/!��.�X�G�	9C?r������EsT��dqRgFm�i�%�]z���Y%��T7�os��F@�a#�qU��e1�u�S��g)\�U�kg�W�}��ey]�Y����5���A���>�g~q���N�J�U0~�� �E���!�_��	�BLu���)�DL%�� �)�{U�pg.�*��:�,��J����iԲg��F���H�a�5�l("�Tǣ�L�$,U�)�~&G�s9��������LHf}��*�')%�ǜ$MnΝЌ�Y��[J%�<� ��b��-Y�:�r�6BB]
Kcb��i$9�ђP�k������-��,kE��:�4�QK���Ik
�p��n+ӰOA�J�V�t]Nue���z���`���3��6��R�j�����ds���C�6�6�{!�Ҝ�%U�V���n�ت.��7�2wvd@��A�P�JZhC�}:��z�FmE�!T�Hk-�S�;�����"}t,-1��+�&�Tl޹4�	��#��C��+�1Zړ��%0�x�c@(��~�p��
�.I FT#X�D�~��B�!(d!�%(]���6��9��𘈜�wY'�P���o�g�K��t�iHc9�@@��3!�l"�8M� ��� )�B��j�t,B�jK���(�!QKM��������	Gtb����ٽil@\Wg\��PH�b�7�a�n��V*C�?D�oy[Q$��:[u�s2�ͤ��}Q�kZG�
s�RU�V���YF'+;/O��DG) ������pI���W�RB�A�9�!k�Yb�W�U�����R��U��1����%.ρ�]򲗾�%7~)�t����6�L\.Ӗ�D&0���gB�Դf2���LeVӖ�7�Mn�s��4�8��M�p��|�4���u�ҝ�ܦ=���x
���?��O^�3�є�>�Pg�Ӟ�B�	шR���\h�d�����(HCj�+[,PG;9����,})%?�RJ���0��@bzӚ⴦��N�ʕMlC��@!��s�Ѧ4�P�ՕVh�I�)V/ЍZI��F]P:�������Ne�S-��j��Mc�S�bխHU)���Ӷ>��x})S�jWJzզ��T�
Wº��~�Zw���
̕�guj�Uv�U��(�f��ұ�5�F�)j�ځ��t�Y8j_�*[�` BPji�*X�&�����lw�������I"�%��2���=�F�6)(U/��mi)A�nlW��=�w���񂗼�=�x�U���׼���#^�jW!�j�z�;���׽���|���ػ���^ o�����9��t(ؿ�|0�����V�~S}���C��#>�4\���X�)�p�S`��C#�pzi4�o�x��p���� ø��0��;d�����>��s��b"S���5�\��"���|.��,� �2i^�D`�\����}sd�|��.v͝��c�zX��A=�s��{Z,z�8P3O�Ԕ կRU�\�RY��
��%+WלY��Y�| �!�C�VΗ��͒����rsR#�S�^ Eo�i�M ��J���-�w�Sw�؂%-��Zh֖���&����SS�֦�����5T�t���6���Dܮ���"E/Z�u�c��T�1�	Ow��u7;����ۗ��w5*�n��[���w5�IFb���&���|����,(@�)Pdb���vx:�y�zF��yDՍЌ�7�c.�܌�L�h�_��5�
Z|#x���;���<�(m���=
j���G$7���h�Z�.�BZ[���AC�̂n�"��9gx� b�kMʺ�J;$��`����&O|47`�LE����*b�Fm���3��Iͣ�4�)
��������pR�aZ��@�'h�X:� �IM=>�EY/��LP^�3W9jF?�}�eM��?+�~"�^�.���)R+j{��������Ȧxx��'ߑ���ݽA�~�3��1��3=���r�v�<�����P��&��u��M��(�klJ��,�)�yH����0]���X]L�����h��2����Յ���W���@�m!e��R�%��-�m��$eQ ���ל�!�-��}����E�N�k���f������G�����)�3�X�����w,G�5l�H��X�``6����C�\O�X�4���	����U�H��H���u���aB*�
��!�U*èC*��(�`RAޙ��b*��!fb n�����u�*��W���"06I���r!��A� XY '2����2���,���Y�3�a����յ����Q� "ы�#.�VT9V�;���"/RZ$�Z�"*�(��Y�]�tT߭
!N!���$^1���#EV�$�	��P��#�"���=�й�C��蝌|��A���p����ɞ�BP���)���AL�L���aI*�ǖ�}��h�ُ��Ѓ��|�N�]�U��E2�]ݘ��@n��y��"+ʢ�|��\�Xz$�5����q5�E/�FN�E�^2W�%Q��(!c*���H6��e<��
۸�4�GB��q)[�����b�(�C��8�`4
`��)0�i�f[xà f�]ݴj~���f�%d�t��吱���5����%q�+-d,Ɇ�`a�%N^�$
�KOM����޺�倨�Yr'�c�@SPf��M�d&C �=p�0���P���	�M��j��lާ~"k^e���kꡈ�f(�[��E'[��+���dY��9|N�.OVpNc��qv���r*KD'A��$�u�q�'��Cj
���̇��(l �� ��]hr��B�ތM`��[�*$`�M�i@��a�\�k�%l�)�����ֽ�Bn�퉃��~ʑ7fo��⹜�ㇶ��Jr��=ޥ�r$�(Y�=�Vf@���x�������I��vj.����$�J�,���G>)��"��葂�D��F��:���d)��n�[:O�aj�0j�0���#�t@����S.�u4�����Pi����t_'�r�A��5Í��(䩵N]����%�j��\���+��P.�������.�������&D⥉���A�蘂A<*���݉��	���:�h	쨩�h��\��:)���g"�l��kJ���*�T B����@n��Ǻ'i��m��"IØ*$oޫ��߼Ꝛ�"���ϖh��+�Id^'�е�L���#�Rr���WT�����G��izX�}v���9��ɝ�B�!N��;1�R��B�FkYhW�.S0���Z|�1�"W�ϲ��GvQ"�k�FHY�!T�btd'�B�-^��f�rE�v��v���h��b�� &�~'�N��
4�0����R�~��R�����z�����j�㴚M��-
��ƥ�e����nC�&�:&)n��]$JMQ�V�c�z���^����dző�J����xF�n��IWh ���Nꔡ ��g�ͮ/\�h�1�1z�pc��fd�m�J^-)�߶N-��Ct��I̤�%����	�����F`C��m� �*O�J�����@	d�^�%�����H�Ij�h�~�ħi�� J<4��C��)����W��z�ͪ��e�+�1�+�c�΂q�¸+��@k�ϐ���&i��h
���]���bP���j�B��B�|��6D��S,��j�(�	#��pj��O6lC��	�G>�&/�6l��d�#��ސ6/&�V�Om֮	T�����j-�'��*��OT,20Ӆ���(�Ub����.S ����3���Psd����@�z����T3�u�'��#�f���
��`����f��f��p�����Ʃ�ZK�z<q(�G�a�d3J��b'4r��2*4�=&
�'�Z�Ad�ܨ�*X��g{���n��T݄FG��,{H��m�I�R��{�@�ȗ��N�P����gD�
b����]S�y0��j.��3V�+螱����� n�P/��-�AFH�*2�ȉ��V�$�PDe>���&*+
��q��2_�Ϣ��<�����I$�B�8�ȶ�N�c�N��@��#'M��
[\3f�3��_@\`S<!`�گg�K��o	��@����`nu����D�sV���b�@�+�����T��X�u�|��L��ZP��d|��<�|9{�u���Z"nr�_�K��tCOg�agy�"GCߌ����c��"~���ns �4� BۀQ'S�ŐX�#�Pq��-ٞ6|��y�P���g<�'�T=�����Ϻb]@�3o����1��s*!�j�4�iL���i�x����c���M7��S�(�8G���9��z b)qz~�]�q����a�!F�S�%�2��Ubw�T�=B} �h�ǊVf��yp*~#~�x��o��3��If�8�2�Tƍjk���8�6�×k�g�o�p���>���Oz^tp-s�xU�&�k83l�EX�$����O��':0�Ԃ�SÏ�b4����0���NO�T2{��#������7|����o�L���G4�+H.b��X9<��&j�+�,�
�+l���ʀ�E� ���XR�Ӑ3(	�z��z�jG���H��Ï�vQ+�I�:&.�^��#�o0�?�E�v��W;���� R�����3�~<��
�$��>-��.n�4`>�K�[�\�;9/�:]�����|��U\<#���R��_Wy�`�#�п��6�"vj� �0�%xL�$���}�gC �&��<����=i�B� zm|�<��v\��=L}�X�Ylx�������C�����f��~1A'nX�<7I[H����OfLseۆ�5;z�e쉘�*��w4/���l'�ۣ4����s��[��U�����u��I/H����D� �rC���c�74,��lt�VB5����u�8;��K{�a���K���?����\���:��/���� �5�*c06�U��s�CI\��C18�1��ˋ�C�@��L�*;JTY�<����>�z'���E��B3���K�#Oxd�d��� �1��A�6��'6��*\q�ܙ�m��_.���(�,Q'@Q���)�Ă��� Ss��s3�3Tt����5Uu�����6Vv������ $��Ws@XX ӷ�8����9��9�q�zz��$�{���Z�|��0]}=�2����2�|���[�\["[�߽j��i{�8w�@��w��=�� �{ȯ`7.���W�b�}�Q�H�"Ip)M&iM��d���/�G�(��S!N�;����r5g�$�1�˝3��Tz���i�v��lX�c���!ֳjGF��v�۸�)C�+.�bƐa
�)�\�	6|qbŋ7�U��\�v��U&!rf� ��V�,[�|=oV�W4�`�B���^�I�Zv޸�*�3}Z�<w���n���yt�7�;S�_�L��4lar���< �v�c�[�-6k��q�F?L}���a�OS���y ��\z.?�Xko������`��.�[�6���� �ñ��,>Վ�nD?�����,��
�^S1��0G�������K0U|��$�*��4KR�"���*���,��R8�����(ထ/%���1��BL�`�
.Y�i8)�b�Z����b�*�a9���N5%N
}ԑ<�(T�H͓�3$�
<ɸ�.B���B��V]5T�I���W��C�Fm%�LW7�5LDv�R�(�<�d�]��fm�,�h�1ŶӬmP OJNl�[c����=��LcP�q��-j[Q�u'Zt�m6uI�G^z�-7����ja�\�8�p��	6�a	�-R0��}7^s�=����O����6��\�
4�crS�x��yb�����]BB�ނݽ�;:�6a$�aN�U5�S���=��Y:��4�2��^�/�y�]V%�[06��V��[�u����ޛo�eI��}��6n�_	`[�D�a��q�ז<��)�n��'�6e����o"�_�3���K�������E�=�n�v�M�a���7�L�Y�1�Ƌk����ӉGgs7/��g�l߾�wl���?�uț���yQ��N5�U����B̗��0���`彊�r�M�_qkK��G�����s ğ����)�b����w���p�k��4(-���!�Ix%w�BauK�T��l%nqW� �hùِ��:O�װQxÁ�1�:���n���c7���v��ɔ�8M��*��\�V�9��/yg������Ѯq><���H3L�{��N�x���b8l����,�c�!�߅JF�����������k�"
#��5��),�=�AÕ���(I���͓M�$3�3cQP| $�(x=��|�a��:�]�u�0�0���p������K�5
�X�&5�}�G����9�a�{���W�9~' ,�	73��#u����$g�J̎�$Z��?0�(~�LG=	F>���C����	20���,�hN�R���{E+;I���m���HIZ�e�2o��
���$�B�2,��8�CO�T<� @��It��gF�(��XTO��vu��֠��!v 0�:�#���+�k�H�$�iC���(�L5rͫ&���"��9��@9�Ϝ�~�Z�)P�v��9 ��q|b��SFe�q3�8���T��i�lҜ*E�nBTy,'.���&��5� ���N|ִ��,T��5��<�ECQ��W:��ta��US�Ƥ��p�˥��ң��$L/濝6���O��k*�:xf,;�<�@�W#�Y�7�*6I7���;b�;Q�.�]2���Dw�6M�y�T�ﶚT�W��#a�9>bN�;~�� :�u�a4������F0���Fw�y=t��芷���f�򸐛�K��
��9��G�I��B��=\n�Z
=�k�8���fU�uK��$S�
��nt"�j1^W�w��o�h�3���\u��C�3�F��\����wLv1���Se]ym�%Ю�0�gt���ٰܶ��+�䐚��$�C�T�ǡ��w�[��ԗv3�'��֒��@k<� �Q<��u��L���N�dm@�Y�h ;&��
ނ^���%���w�i�����6��Zk���ح�jDc���5�cd�͘���6�e� �O�*{Ò��136������gX�]wC�߬�\N�
Wc�����]��Z��i%2*�k[]�ئ�%��I^�Qzڅ���mo�%���
/�(S=S��43���t�D�!6�z01�u�N<ݙ卲��M�O�̝&%���?����\Q����^t:\�Os�cvLgX,�<�ړ�;�dߙq��c�ࡪD�p2�u��a;��c]c��m+[���J��%���v|�L�h�M�y��J�-�q��L�̟�����)Z�����^��
 �����k]b�/��L�6O����`�3�~8t�$��-�otCAW�4��7�싏~!~C�[��p~�t����pJZ�V�9�z,Z\#�&*��8����Y������,zT��I�H/�@��@�mA�TN�:��b*K^�ʲ�<��M~����H��Θ�찶�A��T���.�,�\&\L�9��e��CQ��@����G�ޮ��cO8��g:t ����	؅����L�X�.� ���^�x�,�d�Ic���p�@��"P�mL�:�������o������p"��Jq�&�r����X�+�F<�Hg�c������ڪJBr���	s�)@�޲-`��=���M`e�y��^����e��Z­�tm~�@߰��&�T�i@�by��øeݾ�����P�*���PuKO�PǑ��M��1��8��4��Ϭ���������%ζ����(�,�6F����įb�f���m�CI�I�>�Ep���B��&��Xi ی{�ʳ��腱�e�|g�g��h�ȱP6�
���*Ќ�$k	S�t�i>��tΖ�ϩZR�h��-2�Pn�(0���#�Q+���<��\���P��'  -�cԒ~ԲH� @ �rs*̈͜|�c ���K�t�W̼V��`�����2�Ҏ٠�q�q|�O��r�̒�0�yP��0Q��M�����Z�ن�]�Q҈�
��S\�g�������-5�-�r7�j��-�7-�7<�39Ѳ]��]g���)��Ր+�;��+[�KO:Y�I.�3�2z)-/�l�X��.�"*��g�s]DƘ
^����hؔ/#����hpd�H*��?����C�!G��*��P��NL5��/X�����l��&�4$6�B.�-�瑆��% �j�ޅ9�"�<�r��3G9=�H�4A3I��:�0;�TIKh;9H�,G,��6�k8u�r��R-P}qq�=i�P�����ǚ�cq=˫9:�q.4�o�h�r�c���Ԁ����q����l��Q1#�(���{� ���@w�Kq-�S�Bt���
U8�f��.y�dRH�Ò���o]��ǙUG���� 0f8[d<!�7�S7��Q�:�0J�rI�UY��I?�;��H�5u�0G{�T7=����:!��d�[É��-e,�n�=HA�;3�!�m
2�&j�@�1B�G�xJ���v�A����H{8r1U��HP}H[�(0�O���4�
}[}t]z�Py���:WM5��x�6�rj46cW��Tn�5_zU�S-�9�t*/0WY��g6Y��w+,<�1y�9��~3W����.�1R5����MqOQu�^�>�ß���x���s��ԋ�G�&'���^\��4�s2��z��3)sESb
VĆ�4���-e�F���nEs�;�/�a�(�	6�4-M�W��c��� ������C.QH}�_��-��Z�Tת4.��83��0�<��i���±�L+�h��xCh�U���HA���GgVc��tfX�Pd}�]��[�4�^�!�]Yp`��?��N%*^t�Orc42A�U���_����>���`Ԋ8cR�e��U�/��S��Hd�u�G-@fӨ��C��^hf�dKe_׃���:f�G˓e�W_�sg�3�����xcX����uōJ�f_�,	�6�X��Lg�ɵ����p�O�5��O'3p��>�8O	uF!��uˋV�4nh*�q�P�_�D�arm&3%u��uO�}SC=��g�m�Tv/���*uWW�Jf���֐S8+k�IQ��w��%�Mo��5��3h@��GAf�ؓ��rɢ[��ˎR���l\��C.�5\׊���-�~u>�`��Ю7_����������� ���[��J�(�]��y�ot.����t�hv�;8�ay�1�*7�E#ٜ�a��w�_�b�I��`���iq5s��+��.��K�vR��!�K�t�@�I��k`3�lmiQmE�n۔�$��x ��WP�6�8����6ے6T7 a1$��m��UA,���hq�F4�P����/�v}�9	F�oBlK��WڥQ,�'E�r.��i刞��}R7WK�8�!��Y7s�8��!ՙh��h{��Z�}y�x���Vz%Vv���￬P �V�p3{@�:�� ��	�oL�IXn�"��s�T�P�V;M�P�i���\pW�&�L��Mn��\�R܋*Ơ��@Ž$�S� ��ZNa
\��e;�̀�q䚵Ly)ّך��[x��:�X��:�DG��2�;. -��В��2E�«FG��V�F0�F��2��>/�l?��T�?e/�ú��2�[��#���D�üKd����4کF�8@A���1d.�����F�8���� `˛I���o#mv�˃S#D���3�	l�ļ��L˻Ev���1<)��C§���Ɓ�e�\����ǵÅ|7����bl��3��ٸ�<�axZ\�$�I��ś"�b-�B)��$~�$��"�B"�"��	#vBw���)!�b��\ϓ��a��< �7��w^�(`vl�*����]B ����|�M�ӂ�<��x��P��"������7}�&4}��$%~�(b(���b�]�h��K�̿<5.�˝$�-y��ٓ���Z��U|�3y�ES(�ڇ��M�pe�)X�P��[���+�;Q �=�;W*{�S��c��C����S�  ����P�A�`�A��3\ H�}V�J ~֠
�=4�����A�ܥ��X�]�[��e%�y�)���:��\�[��ې��T��5C�H��_�u���G�Ap��$ԝfZ�~�L$c\��eu�j���64�,H	��]�um�$��]:]�Gݏ�h�+���?��e�����Xg����op�()��<{ۚ��P�i��?��������� 3�/��ԫQ�m)�Ly�n����x���~z
QW/�#�t F5����M*������O qOL���_t�t�2�5̤Y��8f���<�d&zk��/v����j_Q�� w�?A3��ki�%�U����+��_���*y�ǌ��7x+��{~#eT�"?�W��8Nh�ޛ�H��E����� Kg�,q ׉��a�j�7��0�vMӷ����m�ЈB��ZLI�;6Q�+�KD�c*;�Ym/d��erʖ�-ҽn��ӕvsU���7��2�ȧ����"e�GiT����	*:JZjz����������&���)k)
�{X��{�R��<�G��;�L'����qpmѱ�\g��qE͵lP`�Bn�&�%��[P�n|��+�%,���Ⓓ Rd�A^&$2l�.<$�%4�\�r��#�PA.�ݻ�`�2�ҩ��������,�j:���hGBn�ɢ�CO����D�TaV���S,[q�p�D��رd˚=�6�ڵk�F�T�]�Iqm�������Ǽr#D"0�wki��8����5N�
|3v;� b*zH ���ї��Z��3:�@��ή۾�C�4&��݄o 
k��x������2�&U8��T 1�Ⅴ�
�Sj��zdE�1�9�n�w�p�������M3>�aH�u���q2�%_i�]���V�>a�NH�X�UX	޲`X����SV��WO@\UF�U�S2�� C}�0��1�Dט�A}E��9�1#RG���JO�v�@����/�Ǐ9Զb��9�[n%i"~?�4�`6�1���1��A��S;cZדG���p��]0D�tHm����M�{���^j�8У��3�T��QT@0�`S��%$QK�9��6�r�ޑj��
k���Jk��\�Ղ��}����>zbp�-"(	�-q�v�@��M6@B��[_2���h4�\�(FT�U�Sۍ�ƸG`&�ŕDq��[,~Sh4��T���6ڸ�4���+]1��#��o@}���	%��*��	�
���kp��<W�&{���2�Ls�6߬r�$����}�y�/7�D�P�0��H�D�f:�`G����h;֌`���=fH���D�8] 蒍����Gj��<��U4���~��Y rS�	�b4g��aT�tC��N��td�JփgX=E���͙4M���&5�C���� )S�6N����<�}4��*b%$���*e�jpu��\���5��U]>��r'1��}���Xp�z=�q��%���m_�J��;��v�
���)��w-0�"�>�T%;RS��U�r1�\yѺ���dAiW�>�/D�T�ڈ8�upCY_k���� �1��2(���QP]�r��4���AdM�إ�@�TgU^�Vf(�Rlo?�+�����Iq�T����+aHg� ���'=E�(d��Nc���	xV9�=��r��$���4�^��9�xF�<��@
r�,��WĪ%��\ۘ�$*�=�	|�� ����0Q�0�>2�F� ���e�(�j����OB�o���(�W>.�b�W�/	Li1U~�b������T&!���e�6B�a�
|�_��aƬ��5Y�U��V8ω�!AS��d#�9�}m�/q��0��m2���Bо�=~Y\�Y+���zEe�3.���`Jt��(Zx��'�C��7�6���1T����7UήE��G�l�ͥs�Q*¹����X��ꆦ)�@%h|�6!�K��q��,y��ăS�����8���)8M[�dsHQv5j�KYK�8v=�iK8I�D�0+XRz��!\�4*�Mwǳ�]�F˭F�!GzL�"'Lҥ����{���R�z�(e�i��jv��%�\�D��"�d��<�fq�̢_��i���SM{[a:خ�fJ��\ �8:rf�P]�j����M�7�sZ�+���NL	)Ix���oxÚ�r�&W$�m�Wk�{� 
w8yhe-�@�2S���-A���b�����X_cZ"�Y��q8.(� O0 U�`���K�+,�a����v�UG�:A�ۢm&�K�4C��$pρɆ�OW�Ɇk ��ZJ�9�%L��X��
���u��]�|x >!���k��m0L�#��/�(.�[T8�~��w�.hP�g���Spf1�9�
�Hm)
\nH������ X�-3��Of�?���
d7������hT���IP�2�)�J�.&�F���eC�"�d\Hb����6�K�t@nF1�ĥB�X����$G�y�37�#�}:�Ty����E*xYDD
\%����!������ꀄja������)�Nb1�� `��� ar�z�����Ko@�{��^����'^��32�d��	+U9����á*���4��W����HE�1��5��0DLt�͌N���vs��������`�Ų�I���S'H�&ٹv��*LU�X�v\�z�G�1�j��غ����Ҥ�t��J9Ue�恤уP�yRTK; m�OK��6��ȳ����c�a��7ӱ�:3��p�	>�+��^ľ�/�;%hH����6;>���w�:�߁w�ߜ��y_C�W�Q��LK��22��v6ݯ�i�҈E���ևj]���Զ����X3ǟ�y��G�A�tلY�c�K���ǉv�w� ���p�����C�G�6lG��.���lFۍh�t�̗��2���ӭ&��f�"�@o�n�Vz��oEz��y(���� `�3g_}�c�0B�xoxu6w(B7?�qRW|�c�FXs�Q-��l��%g'%��Ej�)�G<�XN�}�8?�T�ZF:�R&(o�J~5d�J`���-����-PVF�0c�Te@�b�Pf#�5����e�xN"A�4�"xn-%�W{Xg�Pdwfy�g�y����g�ho##z�Ɓ��L��X�|d��N���2.�q^�#�A���IbH9�|�g=�-Ʒ�V��Uˇ.��|�}�sAA$*��^�¦ֵN���`�]%�[�s+!�|S�m�w���n�`�@�7��nq�P��!o�D����Ѐ����5�|�+�E�r!.X0��xw�(ubdW({��q:8V��A��#"�HE�v� da�E&;eZAgqg�)+(F4*�TR��c	t@R9U�)�$G�u`�a�ԉ���u�TV5qd>f*[�>n%=���?�{�v;9W7T�@YfCH	y��x �m�xI�U��X!�8	�er֏�fLCyʃ*�&p�����sI��dy�2��K�X�]�mĸ|`}�e�1{>$���9�(��1s�D�ei!% N	��),~ə�t*��ksrB�$ ��)#�_���*�/E��z ]�F�����G�o��n�SY�F	8�&��z����}o����P��mu)��>��y����h��י�&gIq�㐚Y��$�O��u�%��$�鐱�{l��,x����9�G�$A&�G�HH�� I��`@IQIh�#Z��Y(�crE�F�����Pq����`������%��Ɵ����e�pY�x��I��5Z3����HYqiA��|��0�+:)��IB0^+�iS�'5X��8:�j�T/�������.YH�!�v�HYA��k��/�kcP8t�c��R&n8c 5�@c�GC(SmgZ��s!�1�e �j�Rj�	��ҋ�B�0���Q;:�6���
+w��ʢ(���
~�񩥺��W�eb��c���(�����d5`����7:;�4��Z���:%�a�a(����G�R�������I���Z��r����ʭ��~��Z�����J?�Z��
��ڭ�
����]�����̚�����瑯�*� ˯���ʮ��K֭K��Z�ৰ[��*�	+�����ѩ��Q��� �JB�w(�b�`F��'+,;x/�d�^cJI�7�3��F8ϒ�L����C��_h$<��2K����>k�CM;���@;�2�[T˵��Y[D �V۵_���d˴k�Z[�Z+5m�L�"mk�U+�U�1��e{�<��~�]c{�~K��[۬l���`����e�K�`����}븙k�r+��k�'����qw������ѸN˵�빭�����۲�+x_��!P���,^��� ��[�X�,p(W�)[�-k�"���K�0� �뼲;�Lֲ0Pu.k,X�����8G5�+&kG����v��0N�s��Q.�K�{-�{��3���jϻ��[B�k���}&���/��~�U�՛� �Tu8;HVR�������;�|R��K5�*��+���(���"|G�ɻa.,�'���{�8��Ƌ�;����6Lĵ�C��A�����Tb�L��;�G,��żY|G�@�I��_���+�cL�u_���kl�k�(���Z��5?�����a���1��ڬ�ڰ����i�e|�����Zk��Llt����\��4����[��Z��(����ʔ�����[����r�ʯ|���ǭ,�p\ǣ��K�h|�e,����'o�+<
�����7�Xd��E��{GB9�Y���h�{�c{\wIȉ�"�<	چ\'T��EѢN��JdJ_3('GX�q��Uq��R��$��uC��[g�F)-JI�%�H��)'�Y��X�b�5cI9�I�Cb��,(=F���XIik(�yy��E�+��f1>�Z��+|�ry�NP6�7M6��S�s��,lM�A϶i�{�5�&̦c�mC�5�S�@��?�BFrz��B�@����Y�G�C�ֆ��tp�az#�ɗY)�5	�1 ��6�F�Q�l�l�fw���{�{�
��CkʬՉ`Ҋ�mF�~4����Zz�H�	W:_��2}�-�ٟ�
z��'}�4}�W]K�t�vEͽ�s�p#��QS�Pr(�<@9|�ɒ]-JB�W8����Md�or��cۆ�;�m)BYKy#�-���*��������ګ�9R���O�sM҇5+�bo�x��wV���ҏ�Q��������Y�_��D�>C̀��ɜ�?��Զ��z�N�|��^�q#��ۍ�N���7�k���l�6�P�u����x�#�~�U؎ä~J/�����G��~�&�B���z���ٞ0L�R�r�.��������V�t�����H^d�aj
� g'\��0�&�<8r2�ł�T�G`E�"���wjE�' �"zuC'V���_�uӦ�X`��	;�}R_�Xh�#��Q�T�&WΘCtԥ��9#=���y��=���%}D�=�9�=�-G��jhDި�u����G�|��3V��F.O�����^���b�������.����lm�SX�h�kB�F�r�/Hu�բ{ �~e:�Զ� d@���`ّ�+�w�D>�D}-#�Y�Y�������/��1��3:�1�����%&�dG6vw�1b�����Y�P�@�cU�� �^�>�䭃6q?^J�]~�75����0'k���a��a�	}r~R�@�Z�$l��7-RK}��i�ځ>���EX�EV��e�8��:j���})����H�]�d���*�&M�^}�(��p?��*�T��B���մ�پy�m���7�v*�^��cW_x������hO�>�i�>k��Dj�ۗ�������k/�f��+m�5����pzp��=W����t�ꊋ�����a8���Ɍ�^�L2�A]��T8a6�����-�m�Ux�2�P�ʜ�0W���F"G�(�&,ɼ����4����B����0-�6�#�/DKqR��è:�o��{��턯��xD&�Kf���F�Sj�z�f�։���
�_oY�ʄgj'M���h����_�yQ�������(�8����;��ěP8�8H���C���<�9��+,,p��cl�[TD��P�-���Y,��� ��!&��d+:�s�������,��y���������UN�P�}�u�%���9�1��C��t�pL�P� l��r(N"�s3����̠��Yhِ���XS��4Q~���f��(��ܒS�N�=}�T�P)5a�L��(R%p*�������h����*�Y��~Vl�̞E�gl�lǶ��Vn�u�ʭkWl�]h�Z�e�KTp�FH@��B��&7<b��Y��,�^aA�ݹz.-�L����E��V䳊T��6��L�(�3�mqV]L�5�W5Z���G����8�S>A�
�.���Z!�e�ݧ%�t#M`TpE�^�z��ݿ:��#/ɤ1O���I����-�b���!�Ir�{�-�֊�AAH�'7b�c�&���Pl���P��g���̰ȶB��KD.�+p��� z�g� 8|F�#��&����1�4tX1�dظ��)�lJ��S�?���L3�D3M5׼�K(äI<0��/3���QA�zйs����P����,�ZT�m�-=7��H�r�1��L��\�1QӢ���N�n�K5�?E���To���D�Gp��U��G�c!:�	�=�2�ea��MX��U�s�Jp�Zk��VV+��r)�Mu�e�]w�������OJ8�I�,��w	`0��_ �U�0@�~�`��UX�{DaNö|FV�a��$�z):���~�nZ1NY� ��f�%���'���X��?j�$$F��Vm-ޙ��9}���"	b��U�щ���� q8� �.X��!��h%����&���6XE+Z"��,��>x'�p�7S���\��<©I�Ok�ZR�Ė�?�Lϡ-���溱��~���������l���\�XP3���n)vO�|�\��%A�̷��pU��Vbe�n��ݠ�#9�����(��jE���}N���3l:�������}�~��FzW�_��귁���x����F��=q�`%8�|}'p�!�$}�@b������qE`�*a�0Ǵ5��*�^�";Q�ev��n ��W;����Ľ�J�n�;ԑD�*dZ��Vr�|�,���
�X��em��ѡJPd����Jg���H�����n;� զ71�K�4PG�&QЏd ��81����[`����� ��J �@�!�VQ��8���u�����LL�up�!*D;6�%S������n9q}�4"(�>���Y)�R�De�3KP�,Y����2Үlcg�]�t�=[e�2���6AЋ�x�A�t� ��=�[�����$r�nd>��O~6�������E�(�i�A㨶. t�Đ�BQ��a3vs�%���/HhY�eፍ����(0P2-~8V|���\#|��4��'n��f���DǞ��I��[T�,]�;��;U�3%�cZE������OBʞ&i`Oy���ӊ$�"�C�,��;��
-@Eq����bU})G�7��+sD�:ڶ>�s��C$�i�~Vֲ�ݧcgr��:pKԡ�
N7�s�r�����U`�d�����H`
F��)aw��ge�t��L��	*��N6o�KF��}�c�0E�[`�Y�[tL)b�6y	&K�;���f|���d��� ��S��ȩ��J�4���d	-P@ό�J�c�����k,�l����i6)U�c�9Y��0`	�0C��P*upnN#��&I`�7��<�X;'gCbiQ�2f�!��Ɖ*K`Z�"���
꼜��.Q/VT��#���g}Á%L�b���n!�Q���w&p�AіX�1�M����:1��o�s�P.tE��m^��j`Z�B�2��NņLq6,+c��h�xK�s��ʣ%D�U��C�q�2�w�Q�}�+v�4f��R�1�2eyG����\EV"OEz�=�7-�^?�{� �Q7�-�9i�	%��یʓ%s�{f&�9N(��gnw��@q���c�D6V�z�C-��-���1�d����[b�A�߬�H�Df$]�͆&T�t<(�&��RPf	d�Ie� 1eSfl�6
�/�>�Ã��!{�}�tڙ�ޕ�r��3	6��5E�\�Q&m	�7�.6�Vl��P�I5Mjl��F�4:T�-7E���ګ��vֵ��>~��1ʴs�3vԜDz��k���s��YD�Ɏv��6k'f�[���bv�;n6Aݺ�}�H����v��a햘/��x�S�팟���y�L���<��N��s>@6&<����ý�W��]3��G��/��IOx��>5��;�[oz�ۢ��w��_���>�ǖ�g��u�W��R� ��C�-!�PH�q�q�����k�P0�Cկ� �	�_�?�/q!:p~^H5��(������ @|X� ������v������z ?Ux!�p����h�?xp��@��@\��{��dV�@��w��A� ?D�3��|���+ ��Rj��jA���TB��@��%�)DV��'�@~Y�(IA�PT��X?/4���/4�0�?O�C+�$C(��� @��>�0��@ĭ�:>2{�TH�9d��Gl��8��DGDAJ|�J�D���L��N�D�P܅P�D�ELØf:�T�G��S0L`UT~�EM9�X�DS�EL��G�ET��Rt���D�FN�E��KlEe��fFW��kEO'l�EI,Fg<Fm�XC��k��G���`�ilEO�
n��Q���Gv|�H��}��|��~�F~�D3�C����+�P��lk�Atȇd�B�q��S>�3�»H��<ٓ���=ޫ�N�Ƚk���;��;װ�[��ܣ��Tɔ4��s����H����ɝ�I�������I�l���<�x��cʟ켚l��ɠD���=�|��kJ��I�ʳx��\���=F�ʫ<�s<�\���T���˨�����J�>�4���G�s���;�#L�;̘�H��:(�H����|��'�10m�"�q��	��*q�&\#/�x�9��:~�]� X⇏��QK��0)�.�@dD5��
����<��:Z���I�pr��鈭t$���8N輎�h�n�$쀖gB�@��z'�|%ϔ���3?�C��̆���t�	�L�?�L�+��#(�x[!�R5j�lٓ���1��L���X�#(��"�ˠMk�r�ښ���m�O|�'�z����32:"�������<�"X�(�t�=�F�7�xPlp�#.ɚr ��R�2�L�h�Ƽ�	c��d�&M0kS������ �T�߼M�Dl�1�'�QP��K��Jh��[�/}�TSԉ6ooZ-皜���\���>�/A����Z;�ݬ�ҁ���Rd(�6��K�����CEf�S��m � %��*uSF2Ry�>����s�X��|�� 7�47>JR���*�,	90��}'��R:P@H5M�uP����(
� S)R8��8���Эٮ�{�������"��*c�S*�x�\�(Ƀ�(.EW}+U-�(�!�;��׃k�!�
B�j��7Ѿ%�Պ�X���[��Z�����4 S!ԼhӖ�컕IMX�]��H%�M^�5ТЩ��cKM_�5?y-�Y	l����.����ُ�T�=�>(UX�T�h"q'q���}�$�1Xr���5�Y�TU���Du������]��}�Vű�۽=�4��5SR�����'WǑբp�1-V�Ȓ��r��j�$�@��i-�B*��6l��*���Z8���Q/�֎9��r�؝�Z�<�Eկ��ʽ��~=���5��n����	]3]�d�!��΍ω�U6����u�O�-�Wź��]X�R.5ۖ��U�[�+P�1[dE��a�R{�Sc�ڝ@�9Սc�$�EZἌ��ki'�O@��̴C	5층M��1��X��&�=����Q�L���5˘����^��6�.2%+��T�SU_��=��'�|������9�XWE҂\��O`%QE�u�a8p�cՄ�-���g��}���9@֏�Ϝ9ގi��'v ��J�L�\q�P�Z�,6Q:[b������v=��`t4I�����5p�3J����߭�:�[%��0�U<��L��A:O��9��h��`��Z�W!eQ�U�P�՜b-5�ShO�Y;����ىY�]�_��N�	ZS���Tj`�P�j�XJJ�`�����B�5��f�`Z�h;��0�����\:_Ts��������R�M���b�R8��N]N�O��d��XP��f螈�!�0�\�1F�s����}�ZV�8*;HP��q9n���-��u�5�!�2G��m}c@\�m��WI)�.&�6��2F6�Z��яY����Uj#��l*,qch���G�9~-�IfL\\��Ն뱾ፕX�67���R���$4�dd#*�&%*析�_���'�����Ge:%������jeӴ-%`f��O��h#�g�Jdѵ��M�Mfm�K*)��`ټ�f�o±TN�Qa�*��F�ז�z����Uh{Ak�#�����ő�\�e�6n�C�ś:����$�qġ��f6���M]֭8_^���љ�Un��iA>���v��A�������M�"��+&�����x���`Ԙ#�V*Ŧ���ڛ�ّ�*����M�W8ւ���UU���^������?	O�\��^�@���i`�i�>P�{E6��x��i��Y�sA�������]	��
ƷI��~�~g���H��_c�f�Fo%O�����g�nk�؍c>���4����7o���q��i`��Xs���(/��78���Z�pg�S�qg��ʞ�8`o^�+�_�-��a��jl�R����O�m���f�P�⊳7���+S�N���Pg@�^�F@����Qخ���_�n+�Vj�\��j!����	��D��S�vWc�.ׁ�og��d'���29?�� p��m'�7�j]���s�a��i�rV�s;�����c�H�X��:�6n������%q����aWa#s�
I��V��c�T�fk]�PZj��.���6eܸ$ڲ�evmxqO/U;MD���l|CԖ?�sPc���Md� �i��VV�q��/k�����k���N����4x�/I���/$op%M�˽�u-�b��GW.�NwՄ'��gh����p��Zd�ȭ'z���He܈��\5�Ejn/b�nQ�Ƹ��yyyF��nM���ך�ni?]�'���iQ�:���� ������Iw|G,gs�)�V� L��k9R(g���p��jLv�����e��V{�h2�����A�)P����@8&X�J&�~��YX�%��l&|vf�I�����x"`.NIww��a�|���~6��v���l��  ��� 6��KV`��f}�(�B,���{�e{Nh��i:��Asf~1I��	���%K�@]K/e�̝���:Q5�SK�5�%��EM����P������=��h}PVZR�T|du^V:j�N}�����������������������fro��kr�b9"���<[��<X_cgkoO��	l������,1�@1ɠ�~�^��}l�������R�qN��THf11��IPA_��4Sn#7��|�c!ǒ&O�<P@%JlVVZk���"��r�9�u&fr�o@)g� ��!�Q�K�P��oh�0���fVO3��
+v,ٲfϢM�vm%��f#�*�����1|�h�$�2�}�!�3�e���tG#����QQII;-�.ۡ�dr�� ��'0`$\�x�#B��/On�DR�s;Bl���6� ��5�L�i;#Y���|�5�,y�d���"�)�Z's����&��5�I�ACBQ�� �����UZp�>��?��Un���X����+��������s�7M=EM�@<#�u&�'�L�T^���B�D��/�0����c�$�}�$&4D���%(ATJ~F(�Po
���,�%1yt	q�WIL}�N�d��e�i��'#Xᎈfz#�1W%����-LHy(�^@��Ss�iTaM*	Vx��5���4aURZ���b�����i'��蕏�0! ր#ȖN �X!Z"�1@�5]����&�2�ٖXb���ڈKX!\m5^auA�flJB?��8��y��� ����0��\�?��Gu�� Ĳ�'GP%��yF���+��Ž��*pp)~8�i좆�x�K�f�X'
�-Q��Q�k����p�~�q�(R�S�Q�!�5��mOX��*#��`�Ɗ�z���_�G��A"�D�B�)1�j*B�R]��Wc���Wi��)v-u� LXa�.����S�a1Om�\�I�2@Y������M���D��J��P��\�L�tZ�T�����w�< �d75�̤D[���c����������>�㕸5�R.z��<�c8�iT��6��荐b����x�����rԅ�J}�`յ�Fz�դZ���㓿�� �h�O��T�Ͼ���~|�^�@��h�O���� �w?ɏ������h`��h����_ E������ 9�A�p��	�	GBP���
�����M�Ap������@� h(�*�~-�a�D'Zq~�ˢ����/�І�K���g�3�1���;1ԗ�
�p��#��r;��t|�����u` ���t��k9 �#�Cұ~r#J#��8�H�P����G>b�
�R�a��>쓇ô(�HUz撄� )= I�82>w��&m�<&�(��e/[s��R��L$Y H9BS��,��\�LU�q���"��K⃖�#
�9�o����f#%��?*�b��G*o	OfB�&�\%1�i��O��6Ǆ�tZ��Τ#2�h�F�غ�:j�}jA� Շ��ˋ�F��-بƓ�4�*5�I��F�!�x�$M31J�����S��~@�NiIT��� Sj����25�<T�*Uoa5�WB��ZA6R� =�`U�:�c�j�p֨N�!>}�Y��V��u�u��S�V��ծZlR�
���b�*b��X����L]�Rۏ�>5���*`=�ԣnV��� fK�Զ6��T�U�&֨�5m^=C�*�V�,b)�ٟ��nO�J����g:�;QO@�"�������b7���%�U���a�q�r�GgjS�T�Ф.*^����¢'y�9���ԛ��(��ѝ���q�6y������فˈ�3���s���9�st��:!Y�{s��fBm�J]�r�7��b��	H��[@8&N0*^wj�����'�R�2�.MO�ے����=I�a����oL�����1����������{��9�j^sK�6�*v~^�3i���R �@�����5r/��F	��@F1�{^���`�~C�yΡUx�>���Sᤁ��+����G��XD�%�՛F"�l�V�ZӠ�����k;oz�_���l歭9��^��,��y�Hڃw'D���	{[)�Cx����h�~���a���&��<*Ӗ�-�-&@�(wn/�q�F��]��<��ƒ�D0�>�oj�����X�^�q�������9: �o��D/���Dц7��n�Fy�F��ɝE�p��=:�=��d�qQ�{��g�������ӽcS�T} ^�qg���k`��ϐ�M�!![�2�j��z(Ya4�,35���i�Y�`�+Q���;ĸ)1���o�{�ǭ��9���͐���ۋd�RM$��$<��3�
h�+rE�c2�:R2��Fc.Y4#���N�T��V@�#��c�
��D�y��J_nO��`3�C|�o�l�~w�#?\G;�������\�G��Ёn��c�O�w�l�#�-Jy��Ƚ �mW����χ����܅Nw	���J��v��eڑ,6.�=�N���eD����������	+�����	��\r���	 �X��A�-�Ƒ���Dc�\�e&�Hp`[���ʑP��t˶�_UD�Iɢ0M�u��A�
&H�aa��G�<�	�]�N�$�w���`G�E�\�Y����Pt��eú���Ҷ��R�����L�`��TL�=�j!B�W�]�>�|�L���LlG� v�8��ߑ��C
P�������:��a��U��,�o��b"�a �ܕ�t0�q�(b��a)rΛu �^ͽ���~0�:�c0
#/����J��"w�F�0��y��偱e�/��O8 ߼�6��V�ờ����½��G�	��\�M�!)Za���W`�x`é#�HΑ��š@�E�����p���J��#��`kl��,�
����ѣ�����:�D�U�>�4����[��12a��0�dJ�$��I�c��"�,_.�!R����W.L]���¨�b��J��6��)}���ڥ�f�]n��A�]�չ#�����QL�1N�$�I%2E6"M�NO����M^`%N"�Gh��ed��V���dx��� }�]%������ߟ�\�%�Hfn�%[���$IN_I��g�fhr��T�$�1#G`��4��'0���ͺ���8�<�7��� 
.G����#�b�E��M�B$�=f�� ���#$��6�u!�)�P����2��w��tF�>�Η@f���^�/��1��h��|����Dg��fR�*�#�bc2�F��N�U&
d6����4�JL�6��)񦡉gK$�e
g�x%^
�'z�&*�"Y"L�����Th94�b�f�	Q�t�*F��"��F�]Mm�%�%(b&�Qe��-..j&~~�~��Ri��g�� I&�i�ajG>��Y�u��x��KZ��)6���ե�l'�r"������.^�s΄P@К@ �y�
��h�*�	f#t��xƂ��Ϛ0�#4����G܁F�X���8��g* ��T驢j��]�
���@i�a�$�'i
�k"з��kY���G�m�|�J����%`���� `[&�مL����Uv��U~�U��w�V��ҙ!�q%�aKx=�5��P���P4m�z]��+����	��	��^����T@����l��]��������e��v ����B�ސ�+�����æ`,�@��+&r�ᥒR}�䦺)��50)f���g�ƣ��竦���J�ꃔ$��~.c���Ku��PT{��>�h���[o��KZ�E��#���H�ݐ���Љ�N}���Ρ�
*�v��@tݢ�mݲ)���	�`�?P*�(F���i*C��N�3|*�Q�n���g��Rn%�Wh�.r)Z$����@�;�@�֡��iҰ�ȃDF.e��tnC繣8Z#�S.u���(U�$� l;K��(�Ń�,gXe��bFɏ�:��h��&R�ܨhbr+�.)[*��	(^��\&`eRo8i�6���,/j.�Vn�گ�cE.!i���x)�|n->�K����&D@��&�	����|@Ү6��'�n��؎TK���>\�������/�'�h�⮈IA[���/�V�Q�%&$),��}����Q�����R 4<�Dڪ�pt�		�g��+��͙����2��cq�@gB��^���ʼ��L�l	46�ǶD�ve�i��6(oCt,��պ�:I�E�ј�*��:1�� 7_r�C۰����q ��[�|�	��L^�^eZk"�
)��pD_/��ZA"�ڍ O�G"H�LY���N.�*�n�gq1s����|_��o�����2WT��9m�N	����/Gx%͸00��ߜ��$ǔD�R,�K��˞H����k��� ����ȆB9�D�²��^4��A{�63�0�(�sA~lAĮ���ܟc�ޅg��3DN�L�#<qpR�lji�Lk 1H/��]CS�pT$��"Nؐ�?�t7�,�
��H3�T�_���f��=.PO�1;��S���F��en�s�ʨ�Q�L�Ƭk��� �8���樌q*L����ׅ�!��C�fK4�!�e�����!k\�>/#�nP�*Gfb��ti�F�G6��-�A�|����K�2�ò����rC�DX��и�`8Ek7���l�b�r��Bun�vXH�\4���/��8��SP�4��3v9 o�h�e<�),��>�3}#
�c:�c�q��8�����n@W��ʦ
�'�0y�9�%$p����jN{wD@��Hw�Q��K��]�oJπ�me*&O�7;���*�JQ�	�;����/�v�p�-�nsx�[�{s�vq3�^AgC)�:��Q��r�u�3=ă��(��nm_�F��a耏�6��7�Rq���ʶ%��i$�d�K�y��e�|+�$k�A}^$^fc���z��qX=�?j��z���b�lK���#�^�L���,Z��0�x�ڶ�z��0Kn��2��B˞z�P;���u��7A���爀����`�<[B���_��.�
:��^��h{wD:'pZ:��`qr4GWĬ��ִL��Ϸ������F�ۮ{�����t.�fW���0`� �K�xc�� .F�bGk�بʹ��QD�Q+cRSq�.�oӯ��{�^�0/!n[1Z�@���we��K��P^�od���q%�FtGh�:S_	Y �K霈��%������@᷁�ɡo�"���q��a��'_ǋ��Ǻtf�F�q���`�Gfo��ȃ�x�WG�_��do���@9L�26�n;�L�"��t�y8}l���#��9(�,ϭ��텏j~:�����w�}�8D#y�zf&I��f�40DDw)lb�_�z�H����-3~p>{�s�_9*C򴭰k���w�'d��J�3q�	�,����%&ߣ_˓� ��s³qAJX�~�0pbs�͡����HÃ���Dπ��-�vG65�7,T8�?�{���՟d����.M^^�h��o(���Yx�u��5�^�5ކa�w\����$�آ S�ŧȑK�"��"�����%S��9�G��Jr}ÎSB �N �6��P�8�L�$mz)�B3HWlu�8k+>�U�[�`P�$N��T�s�-�8 �x��F��[�q�ip��q����E3���rz�^���X	!#%')+-/1����<�B�HKMOQMRZ=H1RgMeMpeuNmK}im�c[i�]kw��r�1��OqM��[eu}��e���Sa]������Ӊ��w��Q�Y�{�������O�;v��8!�s��n�f�����U㢿��,8Р/^�T�_K�_��9��*��D�:��N�?�e:�hQ�G�&U���&G*:�3�tRh�Ja+��_7��
M��HKV�شO���U����r�{�n�P{�n��m�xu4C! �#@<~�2�Ɠ+��A��,��ۆ&۹U_�|Oo�lz/�l�������'���n��g܆}�;��鿨c�}�v���C�%gw�ݫP��e[��ů��-�zoբ��.ZGy����&���{�7o�,W����+T�
-/��N"	��!�P�	)���Ed����2䎭Z�D�$q@�,�D�X��@:��"+���J��V�D O��@�2S� 
�H�q�\�
�)��E��0�U������m2�
G,�Jъ/Ŭ ��2S�oԱGk�1�������L=���8�b��ޜ�55��s�D��s�PhO�5�DRt�s�0y�Q�KT2G=[ ��&� 5�mv�F���a�C���SRs�W%q�DUU�cG�)�R�/�V�i����i�U�Y��#��n���.Ʌg%��Ak�u_:)d*S�n�)��z��tQ�����0��I�ɣ��	�$Q
�\�Drx��BR���hb�H��z4�i��5����e��-�!vSN��l��[<Ai��n��ڡ�.�裑~ChD�ݖ*}��o��78�:�%������S[���A�Ĝ�Hi��c�Nh������D(�RAY54�թ�"�A8��[9�f�����ؚ��	��p��0��n=�D���ta�<��:l@�8�H-:T�q�w{q����s���6v�i�s�-9��%ij��jD�NZ�驯�zJ�����_~��1B��#8�@x6������8c�ܛ��2�̴	\���ڳ&�i�j��T�V�-�O	�)��@��=0~�K��X��/|���p�'��}\3����Q��|������}mE�IhHpg�"`�6ջNQ�	t!�`C6����0�Z�T@�N�!�E\_�P��p���b�׳�.A�c�#�x=5���mDZw���io{uD��!�%�-�k�@�1M�������e�~c����ʭ�mz["����Af�N�\(� �5���c�G�;(�pxt��Dw�O�2�n�c'[�A�-�R=�
_�!nn����;8p�wz�]1��I�U�xʼc$6$�]*O�r�7�NqJ��3�'�8�jBO���b ��X���!����w�/�원��HF|�k��D�-���� ��.�C�<�ȕx0���\]2K�O����h�V��z�)��˦�&�aP�Xl0C�Н=H)?*�%��H�$�'�3�}�aZTB�����9�f�:�a���W�V�V�����լŕ�L��Ȼ��n�Ĝ���v�)Ԁ�\�`�
@3�J��V�<U��U)U���)	�� e� ��azӚ�wLǅ���X���ez4|m&�b9�Yf�,g	\- X
� +]1���^$�G�Bj[��S����&�J�.���k� G[��A���$k����s��(�Xћ^��W{��&V��ډ~ᖀ�'Q�]�!�����ŧ�m1! hB���-��Y�f��AAn� �iD�
��aI�6�N�=N]`�5�a܊�(Ex
B]�,2�+LV��2�b��#'%�C��ӧ�)���!;��w�7����Uݻ�"��]���<M��W��t�v��<�.�[fe{��/�	���@[Lg̺t��՝*IF-�V���"�z��7��sh!��d�+Q�|���[��Ŗ. �A)�b�+����L�T/�A�/���Z���ԍ����eHd�gd&�7�la[��~o��MՓV�U�H�)`�V!�R^��#C��2�f��5����4����$Q��.ݩ��̡E������$���3L�!������spa�� ��t��z��җ�dÐ���	���4UGS<]���A���:�>���~���l�-*������k�[Ö�5��͏�M��9���P[��p5/�wre���iW�bҳS���\A�mx�@�W%�	.�&Ĥ�]λ@��|�\�^i�4�ҔnB��kA��<�\u�/���R�!�\pyjظ�`� F�N�ɻs��d�4����:����.^�ni���8�2{nf��u�87��Q/��3�=}�;�r��`,��o�%8W��\�=p`���9cI�mFq�i�)8�J���uӸ��})b#��\�(fC���¿����?��CPz����v�#�_/��}�D����1�\�E(J�N�Zn��)�L��R�!0U/y��װ�Y�.�@���m��G�v������vL�f �vʂH8i���d�����®����,�B��D��ڀf��L��D��	��$����K$�� �n~p����w|�:p�{(�,0�$��0��^O�ZM�x`�(j�P�d�o �$Q��������03���Ɓ��03�a`�n,�� h��Ǵ� I��ʴ^`kn���m��&u
��RF�dP��`�VafL��i���B�	���J��~�V� ��.��0����p���VOp�*Pװ����`	������CT�K�1��>gV�U���H�M䢷.���*VdP�|��&��D�4���+(Gp�F��^(��D��˦�@-���v���]��n�d' 5���`#��$Ս���_�s�t�o	t�Pr$3��*���B�MR���W�?PU��ըF���p+9�������6�u���+!0v����LYm��� @ ��*P��ؤa@	�rg-���2	{G�:Ϟ0���� Ԝ�a��0/x ,��"1)�E8�Nj*s&�j�n,�\ dP�	� RK���O��r-Y -�ֲS� ��j�4�M�( /��R~S/�/	4�L�P����9���x�'�p�w��t�6{���l3�;m���7' 6W ^j�)m�(G�bǄ 6�wР����pl@�T��P�p��U�.65��2A���⳵��6S`Ə�>�(�N�jWK@�k�= ԓ̍�j-�k6��<�$/�l���N�<݀<gS-s-��P+�+�0:�4H����P樑�N�2h(7�����B4� Q6���5m�0�R�-m�F|^�6l.��J~��@�����m�,�l�����������tB�D����N��c�b5�j./�-J�,������/8���T�4�.5PK�1��R�s$�695���Q_�9��HuTHY�U�J��+�ƌ��'��S�SF{s-����No<u�F5�D����=�N1�(��>�}J	�,����Z#	��"Ԛ�0��戰� i�� t2�V-�����.��)�
�37ϭdK]i�?c/���lt�^sph7����l�Q˓Xm�8��;�}TV��,]uc9�Z(VֶJ,�Gc#TP�'--�I�p�89U��)@G57%Ub6K�����.�$���JAd��'I�߮��h|�QŦ�ڤ��t�1��B�N��o}�"�`oT�LS��ԋDLgY3����4U�<3�:�k4����
/���e�UڨTp5=v�p�]Rn/��Z�Xk��l��c�,d�U;6r%��ư�s���^�;6�fo�,�(�D�s!�X�K(�3����S�!dZ��^�_!^�V\��|�g_�otjuw*}�m4`�l�\YO_�Us7`lE0^��赫R��¨��vD[m�4�sStX���oKɅVb8>�D�q���x��.vr�~��ǲH�Qj�j��2jֿj�2��d�au8�b�S�3=!�uE�oTG|6�^��VP�^N�@;�4�@�*0Hf1S���Q8��3Bpq� 2��Ǽ�z�V"R�do���}l�C��XN��@�Sy�p% �� T�c�8�S!ל��~���#�qa5*btV���E�2җxꒀ��>{�I�)Bt��t� �W�3��&�N�I�t�&����h%	[��������	Gz�#�c�����4[�t�Ei��)z� ��i|G�}�s���W��s��P��G���]yD�LU]/��q���-�ψ!/�oW3�@�n���~���7��f�6iϤv�l��g�RБ��Ճ����jƤt� 
0l�z����>���a�H�j���V|� g�JNc�i���k�J���}��3=X�^��t8lxW����kO��v���CY�_o�n#E��Fu3���5��.�B���8Sz�Չ�w��g��O���m��gp�|)f@�]|�eJFr&��Vj��%]f�ufe�!_xA\�^fAd�a>&d�%&HƀQ�b"��%�^���Den&]*#e�b$�dH:(��&�I�\Һ��� �Z#8�b�:�;������{c�z+q��_�Y�^�W`�G���eWz��0 e�r+��=�MG��V@d��S��s�Dn�D��, I��o�dL�ʶɁWN���
fdkv�L$e��"U��W�P�CK
�F��Q$@��N
eON�l�3I�d(�"��.4۶OŸ�;���Lj�U�KֻT��?�R�u��]!��X%�m�o�K�ms ��훹�2��X\Q.۲-��w�S�Ĳ#���ë�Edī��3{UFDD���;=�9�9��6^|3�?^�0`<8��<V
1����=8�R�=���B��Ʃc8r#>�C0� ?p�ş�8@�l���C6����|/��<5��7x����EC'���}�9�b<��<<�˧�3J�uc�5�ɗ���Į�=�`�:��`�#���=�Ah�M�CHY�/]�=�=}r!�5Ⰱ��Sf�3����]��TcZ��-¨�"r��̥���SAd��a#f��+���!ֱ�e�ڬ[4�!f����f���٩]�ͺ�;��Q�����"�a�m�ً]ڱ]f��a�zݟ=�G3�Wbe�= {U?}�9�W�9�׼�o�Xo.)�)��pg]�����uM�@����+�K�a��Ƀ����I���J�{��㛮hK�H0>���qP����J��٫�(( ���z{Z��-�Yw��x�}��胫�:��q������)�߱�UE<��P���C�-�)�QW,�KuS�Y�0�*�2J��>oj�*�Z��ࡋ,M%Ju���tk��\����vkX�Ԇ����o���N������^k��*?������9�J��l :���-?*�+3�,wE_|~��p,H�Ti:U�W߳���s�~ָ�Y�-���ʕ,c���$!#�p	���aM����/�a�g��[5UK�����甆��wҨ�#���%�*� �"k��W���8��g)�! ���@�:u�x�Xi�&šlI���¬ ٷ�gt��:^�5�Ȥr�l:�ШtJ�Z�E����Z\��Ty-2_ڻ��I�:��g�����Ek� +[�>�/2� �tq;��s2�xjo6�����{n���}[r�x�v/w[�1���������|����|�fû�>�"~Į�~�{��t��m�ܾ������������׬�����g�� ��x�얻9LduCL��8�(�r��ŋ3j�ȱ��*���Fć��hBb�p2X�L���J4fi$Y�(	�t�"QDE��9É�h@��zjMGD�IQ�0`��p�0ĕ+UJ P$$�5�ڔJ�ػ����yb_�tb���U�5ǁ(����ǐ#K�\@�0�.��*�'V,�a \2��M��Ⱥ��װc˞�ĭ�?�H	Q����*�ѥ������]�f��:�Բ*�"j\�߳��"`���^�/�H��	�ݟ�`Ż���3l����BK0U�@��d�+���_tj�W�&f���8� ��_�%��x˥����a�b��(����������<�%a l��ߌ�x�S��օoA����&�Di䑴��I�-���<�X�]s���/2e0�\����ZRf]T�9r�eFI?�x6�vg���E��֍V��Bq�D锝�D�栄Z��r��LP(�4eUzrhA�\ʓ`��
��>�X��-@C�|�*g����Ҫc)�(���E���䣟N��䮼����FQIR��E�������H��P��nj� �1i�ՖSm�,�'M�"c�$�P������^�@�	��AP����)2Xb��#���túy4�A.�Y�����K�@�@����
�1�ˌl�RAc�L+C�0
2-c��_�W�\n�ߒ��ٖG�(�	�b����О�jK���PS��]_�4��P2Y[�`�-��d�ZZj�z}�+�Tꄕ�ξ���[~��9!��PD������&C64������U�囀���JX�U4��~(�u^�h*zkx��9}Z5.;��ݔ���h����FE����w-oo�jۆZ�k�~��)�Mkl�����G/��];�ڭ�Aox[�Qs;VE,��T�s2�a��Vw2^{����ѐ��3��#BW�G��{O�p�7(��G L� b18�b}
��'��ᘬq
�(A��CZ��V�ҕQFF�C`��" �K��!�ؓ5�(�_b�ǨpDf�����(D%�zK�^אu��9�P�b���'-/�i	�� 7X� ����f@��t�;d����֮~�3^Rp'>O%�J��d
�<Ѐ$� L�(���T�n��9AТ��4`�p��ħ��L�R���Ij�C�HT�����}sigx�=X����C�֬�(�Q��̥.w�X6j����o�=b�ăN{��#�P�c勅՘q7*c�XW��G�x���[Žܧ�O| א�X��D���E�����s�tE�&��A2�r\k��O5�!�i�k�*R�7���b(?�	M�љeC���p�Sڐ�ӂHR�������e������LgJ�&�Ɩ.�e�l�D.Ɛ��#��X����*C>�e8��Fl��({����h�� �.)��\h�V�bP��
�>g����{�U����+�)|l�LgH���'��	V� �����(�U����R!�J_���M@r�ĚZ���Ŭcy��%�����H��S�M�H�d` ��V�ݘj9`��)3�p!�t���fC��N3�4U�\�~����}4��&)Z�9� L���*G�
��z��0)�L��F	���CC���PՀ�ao��j�� �-1Z�����oC�3�oZ�����=�Z4Ķ�]kS{R]4�9�,װ��z�� �fu2L�nMk.,VYEb�϶0kl��ɨkB��*V2U5�oz_V�Q�N�=N�U|UHEìQ-og�Z���d�eHV��
T����T�Z�׺���DE�p1������-0�A�xP��S\��-q�����2�k�J�HJ�6��&Đ�������xV�_�<��b�&������Ac:�7�pY�B��ix�fSko.W�x����g:�O�"�<`�a��^�UXط�6a%=(�-:1~�:b��.A�&��[PX֓����83�i� _�z��x���_���,jί�Z5�a,(��Ll!�� ��+�?v���,S�l�I[����d{ti�"�w}��xg�
�6r���/{a��#6y U�s�.���\r��R�6�2�z�2��N%�ɳ�f�&����"a~^�i�c�#j�&1�,��D���N�M�@�f�w�	���!�z<��wP�����4�#�h�}V���o�*/�;u�qރ�"JWv�kފRC���X55�>���}�S��2�
�qo�q� &q�1cҤ�vA^�����B�]����h����t1�l$�b��RC�R
�NX���o����"����LЂ�\�c~��Wx>ڢ��E>C?�ϊR����{v-�݇��_"�	�������$}�q+rN�sur
�v�}yh8�:�r=�&�dG��z��k�Id����LVt`wt�:m3b��V�SW0�n%�w�I�U
T} }$�I��+�I0gf�rfwI��"�yv�;��GqF�Ȅ% t�x{wD7*�b8�d�h,.5q��i����j�F�7��}z�f
��� �l�R�$�u�5	��WtdA�0�s-uaTcl�D�,R&O��l�{���DC�P��{zԉj{�{��[¦n�%N�8��y�P��Po�Hy'g� ^��Opwm ~���~�p��"?ϥh��x&�dx���fxb�AY%�< ��=�o��W��(Pւ�F]t#=�%5�7�S��.��z*Մ�h��R�^���d	����tX��
����y�P�E'v�hu�vJHv��K��n��AXfA��Z����	���a(K��0����hb/�\(Z��iB)t�}�Eg��Z�p�U^��
s}>ؐ��[��o���oX3�]ݵ��Tm��^`�i\��u4�H0��&��jI7�6]��u5ceU�ϑ� �}L��e	C9co֕�8^�P#k�AY��(@$�a�iA�2Y��YS49�eE(�7i�]�0-wZ���r��>�g�!�Ri�UQi�o�Ah`�f��xt i�/�8KV���FW9�tgf_�b��ɘҴ�	;p��1e<�i���htUw�xRq�E���\Y5i+�3�[x����E���F8�s��AA��@�H���*�e��y����v$A��:�Q��$�t ]a�
J��Q�z�ǟZ� JAʠ ʟڡ�B
�(:�!������2�A4*�'�z�D����*��<�DZ�HI7���y��4�)�HKj�EJ�I
����k��>�	�`�!�-YK��@e�le���Ȧ.TV*0 q�rJ�^��q
[a�yʧ\
�ku��|Z��z��z����
�}��tꨒ�&u��v�J��{���hH�6��������䩆������Jl�Z���r��vꪓzg�Ъ��������}
����� ��:��:�T��
��j��Z���r�{U��Fl��:�z�����:����њ�ݺ�������Z��z���J��Z�֚���mگ���hjdiZ@�L*)���c���$���8 �!8�nJ���&��?kZ�UA��dH�:�9T��kk�+/�0VGkʩ;7�87({�U�8w�&;�%��w6�h!�mʲ��[����\�l ��FkzC�A˴�G����K�IkdF[�o��[k�˦Z{��J�~�]�B7���)5�e���8�Ak�B��%����o���`�;b���˶ԶNk����A��e˴1�����Qk�BH,������S �����Y�G����	z@UZ�;:A#
��H����ä�C��W����?Ȼ>ڻ�{��c����ۤ��Oj�Ы�ϻ�S���;��[�gA�����Gث�d���:Z�J�PJ�H�������k'��y����9N0�;&q]�whֆ�gI5_ϐR��\сN��T�S�Jh`k84���z�k�P|��p�(|�?sٛ�R�'$�w����@����S�]���ZɊ�|�r!lgn)��Bw�>��>숁#0"{��#�Í9#jq8Y���t<�d�[�V����ib,�d�d���'̲��vt����9H�",��u���r��ٝZ�bzT?c.�����bU�r��-��3�bF��U%h��fH��9V;A�K�3�SŚ�dF6 �n��.�.O-�|2�@˵�a��7f�`B�̩]|<h�Y/)�e�Ҍt�ƿD�buc)v���QQ�eV�Ω�85�:|�d� �m�!�x<+1a�vС�^�4���B ��8�M��'��W	|D�P���+��/\�gV��|l���l� ��o�{[�x�og�{
���g�`����;�4MƬ�Ɯٍ
�nmLT��U��t,R�bex��z�6=���xĂH�P�*�Xq)F,����d֥ˢ�X�%�nAF	��@C;L�h4��e�6��9��s�|���ի����5��G��5���Ⱥ�,L0��<-�ʅ��e!�,]B~ǁf�����y� }M�%u�g�֠���j]������B-\��=׵�cMM��:�ډ�(��`LFM�5���Ő��Ű�L�F��ƅ=Ӏ��	K���wϜE�C�ש�-'T�,�d�5�f�-��`����'��;�����,|��"��~qy����B��)*�\- ������'�/�'�,-d�R���c��h5uB=@=|��̣�*�L�tM��lɽR|�zm����{�ͭD�㥩��d��A�W]��C*�,�d���"�</������
�����������䲁�9w��G-�]ņ�;�'��	�n�Vr+Sf� 0��{.�6QVF��>�]a!�nѴ��j�e���llf����/��1=� ��^�7]ݶsE4>P�6n����g�&�����t?0�~�G^'c;�m%�]�݄q�Ȕ��:ǉS�X��Y��&��1PIr�Dv�=��Qv�Q�>f�rw<�[�ȥIu'�8v���w�2��^���.��{=�����L�*��u� ��^ ��(u�2<�=^��@z��ĸ�����I��@���m��l�e)���Mf�%�8Mt����k���=��⑖�������3C^r�8�������j�]!�->{~ܪ�ғ)Ӳ��|�@O�7�yM���Oq��ڝ���s%��N���N�g@ɔ�3@.8S��*��J�����քU*?����/���,��j���r�w�Րhv_�L-�綕��D�~�� ��V��^Z�"�m/�_��|�-���xq_��̵\�%ԍ�q휞��<��H���J:?��q���A?�cܰ���;�e�Ȇb�|�a���s�ޢ�z��BC�;^y�c-��Cpc�.�I�׎2������YW��_�/Zd�ʑ�L���+���Ɍ�<�rBZ٘^�C+?�~.P�n�7~� @��^+���j��F�O/59�u�M��9�_v����V8$�GdR�d6�OhT:�V�ש���5\���D�hc����������S,�*|������<��C�D�E�G�/���KFLF� ��G�P���P�ѳ6SP�6U��;ɴ���L�̖Ж]�`�L��acE�G���=RT��#���T����9[�i��[�h��t��m'��������7�|�}�~��l��=qC�ÇD�zB�Y1�� ��h�+b�H_(�A�aބ�)�`$4��.Q:�<P�%"�($E*Yď(7���I"C
�������iD�U�+�X�e�Q���P�)F�jڊ%�=!R%��o�V�(H�SvI��Xk�awM�a��1��%O�\��e̙�	Q�P�y��<D�����8�Z��ᴁZ�]8BN�᷃O�IC{P] ��])Ӈ�����[F���3|�&��r }�C'0;vΰ�$����噛��~*�8��n2H�|��m1�~]���rG;s,`��C�4��$�X��	%���^�M�ļ�P�T*��0<�1�6��������\�������-F�z��G �r��zLG�vL/	m�ꃒ��*Jl2��m(��I:Xj�,���j�)J4��+;q%%�Ҽ0��������=;؋O��2�S*@���=���);�"�P��iM��,4�G� �28A� P��SOx�=�*0q��,��J;���S1h��?��RN�s<Ŏ�'G�Bc�Hd�UvYf��"<��v%y\���(��)�T�<?r+��l��-Wg[�L��u�8�e�;��Rr�q�X&	�Z��.��j�P�_H�A���Y�OĈGݴ�F�A�	�p�P��x�]rT�@��/vX&�9	!��%�`gs�yg�{r�Ј��Z%������b��W֪��%0��<�4K��:�z�'�.��si]!W�8JK@�DX������
��8���Y�jŕ�� /L}��2�(cJ�T\"8M�֧RN��ֺt;#5�#Zc�(q� �Re]}R-� Tօ����`�b�""��ׂ��ͿV3K�V~uj!��	'᝙ZX�� �g���{���՞�|!>��dsM�	��ڕ��e8�r=��®q`0�+�t����E5c
uTA5�	�A\J��y�:t� naz�PB4��~�� ;aOt����'�Ғ@f#�6,���gI.@;T&;�H�bRH��� �:~�;�#����Š��
�P,���mQ@�#���wF4�Q�:���t3	�'S�iЄP����u�#
�
5(:��$[��dҥ���@c� �Z%����C �����ln��H��N/�xc5L���*��&�D�K�HI.ׇVD$ny�]�&p �D.�����L;:������>t\��'��T�ƕ�8Sr�#�*�d����5"��fw)/��mL��8�5�S���dd������B@������K���9!��= ��еq�$�3D#�E.�ㆃJ�&�1�v���HV�|�{`�"�$>e@����#��/�A�k�s��a&�5E�<:=$p,O�ѷ�`S���kY�Ҳu�H	�V>���z�U�c%뽠 ��]���^?u5R��UU3Q�H�Ч"�p`�Ҟ�����E�B��^���ȴ$'��2��TP�_vR��H�0�ͽ�@{��h��p%�S5=	K�!&�p�%g�����n]�i	�j��6�.+�G�@�ȏ�*�T��]&�����BU6��Q����f�И���L��]��7�
�����]0���+�k��>D~�"b40yQy]�k�s�!��%��᷑�K[��/v)@$[���K�V�A�)�,k��V�-�LB��~�s;���.�n؉3.<����I�T��� �L�a��P���:���e;�f�\��'�m�0��`�E��e�����K�Co���eZ�4��0��̥�vf>
+p�˘$C�7\��4gk�rpk6�����5��Ϧ�&�}��zІ�]�}
H#Z҉>��ohI/�͏�t��|��Z�h^3�iO��1!s��5R��Iv�5�Y�&@�zҏ&��+�fCW:�d���}ld'K��'���F[jg�4��BN[���9� ���՞����	�,�F��mi���n�O���n�!�J����
�0��3m<	<��V!�o�������,��om�;��.�	����A���F��3����\�����[.��Ǡ���ʥ�o��|�Kf�S��.?�*�>�׸J7w���f �Q�צN"�R��+���@����5�X�����3<"3?�ɹm�j�]L�6ួ�}�0�{�{߯e�q�\�o��Bnxė��t�ÿߔ���~���t:>��V��-��·��|���#���o���/O��Q��ݯ���3����Y��?b�C_z���O꼻`����{[�w}�/z�����=��3�������|�_���J�~�_Qڑ|�O~�{�Ou���/ד��SN?��z���~��C9D<L�(X6�k@46�b��[��`�5_�776��5B�4E{�DӵS��( G@�<�FHAC83E�5D��TA<�t�>���M{��1J(�A#|�D�7#��3�%@BWXB4$TB�B,|����"��P��d41L�1�A2<C-�B%<O��gX5�A[35_�Þ��/<3�5@�C=BUs�Q�4^���@��	��|@I�ľ�@�X+�j��ȻY/?1�a
��(����!�T �8{�+�y���@B0�*�<	��j.��V\� z!
��4��ܑ
c�3�2��%Ut(Q���)d��c
��Қ�R����9򋃛(p����Bkȡ�+Cv�7�DJ�G{�2K�L��,�N�'���p��*�X��һX�ŋ��		C-�!�Ō!��
�Bju�H�����J���r�
�pH���E��I 2���+ ���z�m|��������0��ȳJ+�B�q���/� ����S���b��0���G�˰�IU�J����*�
p+��R��κY��1y��� �60W�X�,�r t|�p:��jښ����ॹ�Fd��q쬶� Њ%�iG
8�d̚n���LbTG�"��Դ�20W� �D����Թ�ǜF�)�ѱ�k�S�KPH�J�%S�l�ѩ.nT��4ˀq'��J��J��N���D)!.k+:H�,���S��2�,�{(?h�陗(�,�@�eX���0��wL���$13I7@�� ��LK�����+p�h���*)���d��� �MMG�ɭ"�Q�)*�0kJ�N�Y�I�Q�I�rϳK�������Q�E�����J�TA�ʱF�JN��� X]����e�7���0�N�O�1'�� �:)���p���pCZE�d�A�͘:S�XL�<5��&��Ô̾,����4->�FZ��v<S5iR�����t<�Lt#�,��TIU��*��J}��q��O%���̆���ї�̊'���P�3L!uZ��a���JMl��LO2kQ#�Η�7m.���NzyOJ���j!��@�)Ը�{Q�-3}K-�WE/�TqW���N���2��<&@��:�aD��M��%,�|+� �m�
D�I^������y�ݛ���4N�	�A3��_D�����҇�M>��՜M��,ҩF��T=YWlS,�k��tTU��Eݪs=/��Tr�Y�%�J�Q�QM�Pm�o Z�0� �S��lHudCe�C�-M�VL�k��� ���$u�AL`� g=J#�Qw�"�\[��oh[��Pd]�–Mլ!�kY	�[�qR`HH�hۙ�2�UK��ԝ�\��sm�v�*uus��!�XXBE�%3�Wr$��!JZ��G�{��D�*Q{���Z���<%,1M����9=�Ql���Қ��r��U	ͺ��=-|I��,ǕR��4����e9]��� T�؋5�}S�eF*���=�� @��-��YT��u��@�]ieԛUP�����_����z�g]��%��G���򬰩�'�7�3(�[
>ܫG [�b[OXH�z˜�!��
.a\������oe��ؤ��
?ö�ʴ)����V�P���a��.�\��4��Ǫҏ���4�u-^|-;8a+�	��0�T�S��)��+���B�޿�^ӹb4Nc�`S�@��#�S�}a��@�������_�R���dBއ~܁-�.A�cyS���d�̤��/��c�z��4���G�8����G]�0E�LaV����3X���L<ڽݏM�r�e,`�ߥz�Pe�vŇ��խ�V>�c��a����a2(dj��]�����[J��ǚ۪�'̔99�9��O���FY�^z�XpB�+B:_g�8��,�ܘK۵LK�'��e_���%�S�-$�]2.Q���R����@ig�6��5�S��S:%Y6F-��U�n��p�%R���h�b�0����`!b�Gȵf��iR����mv�F��fF�X���@��h�-�f_~�O�)�h�c.�[�[�䂑�ne�9�L�De}�Y.�!x��r�� ñA�*(#�
�*�U�V˘l�rJ�JՈ��%&��!��i�N�~l�^e���!d3Ⱚ��!�f
(�B�+]ة�5<�UBUM����l�%-R���Ì%:%����H�/NT�m0��mƱ*dt�<Ҋ��n�XQ�͒%߃5Qxv���Ц�a5�.��c�vh� ��V�:Fn�Z&"%n�^��Wg��G��t�l��o��`hbi���-�> �
K�i����O�3)qK� ��Y�œ�M���;�����Z���}1�� l*(�����p�vdY�O�y&���*V����e�������-����O��&���.f��!�b��^Q�yq�i��oE�o)���ʵl��˾.��&�ޔ�B�υhw]�@�>y�s~g?_���+=P$~f�*���Z�д���+-P�<��ME����Q��.;P&Dj��b.e�k�#(
U��j�Ng�XI5�h(����-P'��[��l�tV	�u"��b�tJ7�I�@�ߔ��?Rl,�f?��)�j��(ol-�g5r����qW���R��������ga���X�[����L���nk"��)'_&�Wf�X����,�Gr���e�[�qh'��n��+�qႁ'(��ֺŪ,Z����V�&���xp`b��b[V���������-�u߭���R�X�:��]8�׭n�m�;�B���^o�H�L�˽�%�?2W��qW
M�9����M�2X���$�Tr9nnpZ�"���:'?��S��$��w�yx�\���V'�R��A���x�~����yß�C6`�?v�ƶ�oq7�F9	诬�]#�l
/��v���F��_���7WP�F�$�v�uXn�zi`���������UK��PN���!��q����0
�������a[���v�^f��w_��ƽĎ����ȍǛ����k0�I��9�� D@iм��B����#s�hg�m�{ R$�Vg��Mv �Q� zc�������W�[!�Ғ�X��'��H��'1\+[5]%�Pjh�`g��PV��T͎?*0:��Q�ŀ�������X�#[P�!�V�Fd��昀ϛd���]("c���a�ޏd��,�o�/oJ�����1�i��/�3t��4u��5v��6w��7x���7�pr�3�9Rz6GA��<}�}��V/%W1���Q��w�p�*��"�L �,@b��&������D2�3gy�8�%#_�F�TS�I7�=k	-c�50�d�x��Mc�6.�Vf�@}Ţ�"q��L�I�É��A�`sw��Y`%jJ]4�ؘw���Z1��tal�̥��0t��FI�0����3n��1���|Z���å�����3�П�.�9P�@��^m��j֯?�~��s�ـv��M[��й)�����m�z����i/W=��u��q7?�z��sw~�|p������������x����?��m���p��G�z�շ�`��ÔdJ8!�Zx!��QVa�Ax�mMTr�����'��� ,�8�N$�8�IB�4�8��:�8I&���f4��#�%�� ���8�b�4:�"
RV`H�����R��d�5�I�BQ噁|�{��Z�h�8egB��W7�(#��X���Y��v2�g�fv�$��mIe��৛%�g�u��
3���E4f�'�z�!y�h�L�g�V�h�����㮗�9i������럄>�h�eY�*�.ڠ'���Z�}�e�e�-��;.��z�!5�"�m��	C��~@i��Hƽ�����Yڒo�B�;�<��/�	�p��4|��� H�lq�CH|qġһ��d�\o "S<��<��-K�Z�������+��,�l1�;��2�8�;��<{���-����I�r�7b|4�H��-]q��R���N_��Z�[��)�k�E{�6�Mg�q�p����Ov�y��)�[�E�����+�8�;>�� &X2�l���.$���Xr��#�c�m���IW~Jk����������'%iБ"�9��_V2	�'��b���!-�^N�;�GX۬��>�$��n:��/;1�_og���~"���_���[�"����(������Z�_�/޳?����<���ҡixyJ���;��/V�[��a��E�C9��;��r��$G�砶��~����sB�|�;'4΀�#���P95��DC�'>�i������15�bub3D&��i����Jх�YO�h�������Mx0��f<c��"�P;�a�sR�D16�r&a4B��=�~T�K8B%UЎ�І%��ȩ$��*�>`3�ɹ,I���$�l�|E�|Y��N������V}��`�qXRND�DH���Y6��1'�_Nd��L*���D��|���<�cLae*s9JL��)=�&I��dÂ����.�����|'<+Hu�"4�3Q9�S�b�F�fJ��91���d+�`�A��]���EF⟃H�E��xAᛄاC��ˉ�3�|I椌�&Si.j;�4 �(Ls�|4����JQ��4a�irБ��E��iFs�QJa�Iٲb��3�AM�B9�Ϟ��#��O����k.��lk>]Ϲҵ�v��<����Y���F"KL�l���JH*�bJ��(�\Y�}D�� �8=M�l��TF	I��2��|dB�p�p�2�~ eZ��Jq��ڌ$Sy�L�P�2���}>CM%���5�+7�Ҍ��S/d�K#�b�u.Ü���]����r7��U':����e���2fSk�R����^��B��H�u��}hn{���~wC�����W�i�*X�Y*�vhE������dKo����Ԫ���$�c�M���@#��!XD�H�=@l�(�$�izEI֨>%,!ͬK�p�4�2U�0�{A�N7���.w�,�)��ʝ.��ڍ�~�!�}f7I(�Eꢒ���6 �\��Y�nn3�dY�2�`M	+	���@���R@��;����X&lq<Y	�����-2��hz��ɉ��Z��?C�����/��Z�nR��-���<^�R�ծ~u�u�j��u��/�u�^�*���$ �P�����K���R���8���y��§ tizR�gW�ٖ��JB�w��>�]֣&[�+^��u*:�n�ٿ���io[;��ާP�Z�w���lE����09��eK֯f3�3��G���T�!��j[k²��S._37����7g:�ʦ�.�L��.5�Q��!Ó9���dP5N��.��҅�m+"F����"�zJD����2�)z�c>ѡ?7맖x�)^u��}�8��.wS'�օl���`��W�9Gqz!��d���(��|`#pē��<n�����W��mo"��Ҟ;�	q��q�/���������ǘ�<�%� ϼ��Mi�%�u�b�]��U}���y��L�#^i��d�$�;��/}�v��N;"�b��ۑaN�7*l���yUṣ c�v��pt����}��!魩���+<�o�>ayD��V�ł.y�T@KH��cy��Cq0���c���9�.E�؅S{A�.�����ĥ��� 
N����=�e�O�ھ��u����1��5^Q�������K.P����]@T �I��<�B<$��1�,��ν��u��A�շu^�1F\�A��E O��U���lTR��[<��Mۿ%�X�aTM`��<�@�V����y@u���|M@��^�ޕ�e�g��&n┭ະ`_a��{yY�����̹B��$a�*VK�C�����Q��V,� �}.ޟ0!�%`���yZ�	R>�J�� ,6�%��EZ6`[<`3�" j]�Y�*c#q�c�as5c �3Iۑ�Wu��q"=�#'Z��0�;¢�A�)"�ZW!��������[p�pQm�bB�E^$F�CV����1���0�����e�J�$K��K�Q��@;8�|@���P;��;�#�;�#P%�Y�h��N����`]]�4NAML����YlTf0��r`�0�D��K�%Yڃ�Q\� 4\&3:�Qh%ݙBY֥]�%^�_9ΤBJ�ߕH~P���ݕ 
%b&&�M�Y��)؛�Sd&Qh����[���B��'�@?�f�bK�a���-�|^?�fA� �_����.�X�c�o��ZZ��*C?ЅX(�����!,)�N�R�[�E��@hVf�z���ă��9b�M�]-,$�ş;�%��(*&}�gv�U=�"�!%5y�ҹQXZ'A�\:�]�LhL�/$��Ze�Jb��N(K<�RdT�a(a!�_YU�~�ez�(K����2� �B�J� �(�bE��MLh(��X(/$!�������� >��Rh?�hV�hw����؂>�3��)�_�.CV\�U<Hh�L�$�"��)�d�)XAUxe�Fr�ޙ�����(�J()�Z��$j�FlUNR�a�aڧ�*<y"a]b�'vuؽ'��a��AZ{^�%䙊�,l� 'G�[Eڜ���o�d����*!����d���*�
�B-Bpb n��\'#<'}��'h}��hR�x���V��i�zf�B"�j��z�f:��ߌq>�W���4"*����(�*Q:�w�|��2"/`%�EҮ�k�E)%�Z6�Ur�2h��C��ܯ �-��&_�f��R� Ģ��Qc#�^�1Õ�����2��ƅ�B%+2��jF4���j�lr��x��t��6BV�ES},�f���إ5� ���V���u ���7��Q��V��&�:�:�<B�ΤT&�^�*x@h�U�ls�m#<k����v)���?-l�.g.A�a`n��n�޴��h�%+܊�*":B*n���rZ����d{rU�~ ����m'�*`vQ�F��	�j��.|�7u��+Ej��E`���FcÙ��'�d%n->]-��d-���(�U�*�iR�b���\fȴ���k1�l�l|!�̡K�MDrыȭAmD�Ē��>�H�����ЙD�"��z/vf�3�f�Ri�A��*��F��"DK\�$���I��fK�ƥ��+�%��:囎/�*��؉,Sd�в���:ɣ	/�0��뒕� �c��¼F�*$A^g�".�����y]��>���v@�Z���pAՠ��pu�o�vF԰d��F�@�biz�>�ڶn��^�"�k����J����@��nغ�U��K�&��#`��2������qw.�T��T0��e��	p���
��X�.uz&𝂤�+���"W��2+3F����Q퓉�r}��!E�d�>\EP�_�	qV�)��/���ne��E(R0n 	S ���h��m3X��摦^�P�N��h����Y&{�Ql�b��r3���b*Z l���=w/V-��b�l]��VAZh�D��5��f���X�A�&�L,-(g��� ���ĩ�Ԃ�O��H�t�im�2`}2?��d��T��{�|�^#2���Zo��-�J�tC�᪆+I�TA�!�u�v�˂�t�T5�H��'�pB�z�a.C~�'C� ��uVk�����5"�`�D8uJb��Ҵ�j���[q�*��`6[�vجw���Hz��k��|�xIQ-���dGv)��Pe��IY6i�h�t�li'�u�v{TQk�2��lOvhS�g�g��?��mo��~��,6k �%��
a7�sk��K��T��\��$��JՐĐM�Č���X��|w�,�yw�؜���ب��tiP�ڬ�{��ٰ�͸M�ȍ��w�8���"�����w��|���ب��̌7K���w}���w��͘��O��0�@L�+�}s��)}����7��7�8��hN��`w�t�t�H=���W��,��Ȉ�H��I��� �����dU����)��0��`��@9��O��M�hɖ��`zO��9�8Ux�����ISe��d7��y�o�SO�89�N�#`� z��O�HO���o���O�����4z���9�Ϙ+:���\���ϤYBŗw��s� ���3ӫ���z������?7�6UGbK؁4�T�m��p_6��
a�f3�d��9�k�v���6�w�c/B^�{�g�oo�l�{k �ͦ�e���c;�(�KN����yv�w�#��ѯ�`#�,_�~��5��J��[��8� �jH�}���*N靘�"ڒ�N�[*�p!*�Z� +f�ҭ��R���)�Ư��p�1DVf4V�(Nq��2���)�*Z�3<HǣԆ��?==f-J_�_��� �0�Z�Q��o���uM��[�@F��ZCU[Cg0��Y��o�ȟ��k�W*A�b]�$���᭽�n��ýP�X߳iO�b��	�d�,��X�q���ļ��!���9>S�5�_W�Q꣹�+ԟ�	{ӿk�']��W�q���v��k�3� z �΢���m��Es���l��[�|���{3���*nس#Oj��3�$����9�/5!E�Y�k FE�V�(	Xt�>շ������ �:�I�az-(��A�- ��
a-�V��j���L9Q�Zmk���T���h�$Z��E�	gŌs��E�S�:}i!�-�4y�� �"BʉX�W�ez݄�`�O�0��lE�/�)�#G�(fmb.*�Np�FHl̮��b��Ԕ���t��EU���vԣ7Ww����8Xx����9Yy��cx5V:7'v6���P��2�;�ܔeO������%fk���9ݕU���v�~�Qv���0��Ŏ.�����W�vj�e��VF�q�W�,��Ffzg��S�1�aP�Jo�}3)�̓�H|8�$KrAc	��s`R�K�6u�jT�����h��Ҳ�B��ۇ�@P� p��K��_�y�B��YN�^9�-N���	�W�x��2�ߛ;P�\�th��<=B��'`�'�G4����N��$ I&r�hŒk�t��EA�1�t�wG��MBLB���E!K��J�g�*�R.�l�ȮѭM�Uujv�۹w��<NaմV	��1� *�~|���ק?Q�ۖ�W�Hz�t"�7�ڣ�����0+Rr��}����
-��)�g��D;e��`Xh�]���
S6�e=�Z���p���M
�eP�`�Co:h�Л����<�$�\��J��]�*ϺZ�"l��,���&�$��Ҡ�K}n��ϨH�A���ƒ�׼\M�+�ܓ�=9BN.оR�@>���)���t�$��s/B���D0�4�Hp젓��8�30#s�!
�:ψA��Xe���Z��UUIJ	J���*������ j�au�	?3��r�[���ix�ǡ$4f�p�vG|�2o%igi�Ū�I\H0J�t����{�C�E 
��b�C際~bhXr���Hx5�[�]�Z�Uh����-��p�(�t��l�sN�8�ē� ��N]66JK>�M�b���p�Q[�ޞ>b�e�ڽ�Lk�1T�7̸(��{�
�1���g���z]C��7O��r����z9�J�����Ր��8��ޛo&���aV���}&�O]��΂���$��2WA|F�93zQ���b\�@���p���{����� �������)� ��*����� ΥwW�\n����_��A^U��y^P�j����[YP���k�Y	�e1��5NvgV�
��?9��(�w��"jA>{�0wJ���#���]$���恅s�S�Jƽ���g`K��@�,��a1��wA:�-u�镐HW<�5�y1��i��A�yޯ�g)���G��U:���YN�A�@9���LxS�td<�ZII�s/�M�`�H�;VW��Ў l�F
��*/�"���L�W`t��hb�֑X���T<#ƫ��T�")�	�nȓ�f�s\� '�$2y'4�PrbN0i t��$*��
`~u�MJyW����d+/��K�����F��2�Q }1�!�����	�����?�=����"\�g>�5��pPY1�W(:<0�\'~�[~ ��$&A��Hs*c�[��9�e*o'OF��Wk;9�N��pJ@�d�$ɯF^��菸=���:H�N&5��V�R`(m��x�K��B�.E�KC'/�Ȕ1� MZ�VntfD#��1�my$��
��}�:Scʏ ��M���w-)	 �'%�J{J���T����Nsi���m<�+>�VսҏU����-Co� ��`	[��>�UE�V͡������-e�J*�3��lP�S����%(=����t%/aΝl��cM=-#6�d��|�v+�xꫩL`C)H��e�,Ӳʅ�͌g�g'��P
�E+.m�˖ϳ��D;�΂���٧S����-�f�y����U.�a��_�ڊ�r�az���:�G���IQq�Z�c���Za:WӖ�)���j�Qt��j{P�5ء�X��\-^�S�f����ơV��ش�]_4U�DV��4�Uw��G* ���ʂ8�`Bc|d�^�"ym�w��'Ro��GSQ����i�V�V8Q(����	�)Y�L�%"onWI���V�Ѽ���#M]Z��ݮE�{8� ٘`���@���=ec�	��q7��.�|l�ʢK�@pY�jW��t���AY���Q�u�<K������͋�h$�\lc{r~,`sxF0#x�&!�+7�g8���bM�jh'��۾p����9B��櫺M�⽾���f��f��u�4ދ���������+��&�����{�oi�;�`��_=�Xd_�w61��6�	�Z7��ep
��Kåg�kEsVmēv�\]A�֠i��,]k6NOX��v��������%ӈ�́���--�9�F�i�0r���`3�
��WGZI����h��4��~sవ���s���:�D���2��޲��
$��Q���L�W��o����/mVYlK�X�M���ّ>]�2Y�]e�V������mZ��x3�h S�n�:�C}�aL\p�;�4�1DJ��J<%�Yu �%-�m�CzM����>���3��h�����:��z+��z'�l�_ez�4�4i��Y�V���'��%O��� 1.��c�(�WĄ��@���H �(��	��k�&0����j��"м��Z�K	��.0~�~3�ıM��	@��0I���D�J:Ml$| ����K�� F�@��@m�R�D��S�N)�iET��p0���bƠ���4�ۀp۩��3�d�rnS��Z�9���p�I�����, �Pό��_���Q�h�mk� �s1����#Q'�D�)-�.���3�E1E���SQKqU1��3���ڸ� ��U1]�[�1�o�wQ7��i���_Q1������r�d��3��
G�($��+�cN
ґ�jf��"Jd��1���&�Ց�q` 0���/��d� �1 /i!���A�
r'�l1 � �"�Q!�Q#;23� ��"��J�$3�W�#R$cR`6�7�!R&٨�TR'�n� �(&gq+�$��h2$a�"��%_�"�R(R w�'ER s��� �q��#]�!�Hj� c�&_ �R%� �q�R�*�����r'3�/���(��,2@����U�Q1���WR�,#�֨,e���2Ϡ�43��<39S43�3�",4��;3�b3�3݄473	�6o75d3�Ҕh�7Ys438�33iC8I�5��8�2��:g��f�.%7��O�S4��:�s9YS6}S�S;�S:��<Oc3�f;��<�s83�;W�;Ѣ2�r$S!�$B��1�@��I��J���=qթA_Q��34�nqCu�9�A4�D5TBMt�D8�W-CQ�Ds&Fqg�F=�D;TGG>���BQAeQ�`qD�t�IA��DGtotG�tJs�DAQJ�TK��A�qI{H�I�QL5Q�4Hyq�A��lH�,@�N�b▭�/1ǃ�j��E� ��$�����Q7��p-�d�L�����ë�c��E�S3%�t�8&W�xb�D�Y���US�����??���Vk�V�����k��2
�tp �Xpc�eE����4:�-J��8�����z&��P�D��N�*4�-	��Dq�:`Z�.�0h���~ؕZ�.YChbM���(C�T����LhP��R/W[��la�;t�3b&/���%��q�B(��x#���Y}J%��W���TU���d�(�.e'5e���Bj׉U�Т*�z�ҾLTYc%FwJu_�U�E�H,Y\5ET�a7v��Oa�Vj#"بN����`���A�P��F���נ�eO �UYe�����,(4��lʶX�ne)��Nh�gY-�d��0�@�k�nm'�p�~�i�R�[���؋N�p��^�v���X��K���t�b��tO����a�i�Ftjv���l֍ve��n�pζ
�)j�>b�Qk�jE�d�����
̮�S3�C�vK6c!Ug�j"zvDU{kl`T�hY�(\F�U�OYwV7u��t�`�dW��W/����l�f��G���(wN�(V^��B�6p�q�U��7qq�Uy9�jʠy-�R�w��g��u�5�������ZOhh1�� O| �~T.mWPWEW~���a��i	�tU�ݺ��@�z��dw�j3��7U��
x#/1��@�Wz�XR��ǘ7�wi�|���&�r�y�Ll�C*{�x{�7z�V��Lx��Vuq��x����Ws؏ku@�7U������~��5e>-~ƶ�*�nx{D�R��e� .Y2yw/�B�n����f>lٵ�w�3�
�R�XWy225;�4So��w������	��y��ˋ��C.-y��YL�8/2�{��OD`e8t�nh���؛�Nc5U�8w��ކ��f�i�/$Ǧ�We���w¥��؊�J�� F���l�se��o��Ϙ��8�-���jPS&��%�V}�lf��x�wt������}�~mx��~��ل�|���i�G�Yx^y�5�5���.�"ŁA���Y�!x�$h�F�Yyoe��8PO���N��5�?rgIN�����壦#r�_�Y��9�,zt	�^YdJZ�s��t�����Lb��g��XG&��5�Z��U��_������_׆f�OR�P��A���o���c_�YT{��7!�yB�ک*��č�O��E��Z�Z�����皶0�U�^H��Y	����Z�q��� �#��;ה�9/�}z�������&����Q �<��������h����9��K2B\+��;�	����W�L����:��U ���>٨�U�p-�:��`��q[��uk��0�W7��Z}��v���vwĈ{��[��s�MY�m��M1[4��x}Q��$�.$ ���#6e� q����e,u�ȳ[�b�Y��ȝ���㢣�e@�z��Apj3\�AZV)<�\���,������W��/~�@���w��<p�K覱��D���nG�k��	���D�~+�%!D�V��C���Fވ�M�Ɨ�><4����輴-�ڰ��/2�~����X���K�EX�^����r��0�M�kwWkpďt\�Z�����˭6��\�Ϭ�����ja��v�Cg{ͮ�j�����K�����pG�ҙ�������b�±���L��h��&Ū/�C�F��P�"I[K��F`��ò]�JR��h�c��T�������.�|}�}8ه��t � �|����A��e��A�"�B�ڹ�2I�����E]�м��5����vWHJ�މ��F^�k� 2�k�^��k���-�ѹ;?03��g�� �յ�dv����������a�^T�_�4o߂� 2������F��7�k�A#M.ݻ�.�@�%�]#�/�4����G�
��6��ʘ/�4/���m���P璃�C)�U��+��G������\���+��*ʢ��́ڗ�H���*� 8L��� �E�tL�~����\j��*�JƬ��[{�-$�3\�Ὧ|�F������|_u�-mυ�$ڗ�_Fލ�W;iɷm[�Q_�˙��ñ��<�Y:�>m4���`���Y\ed�5�Ӱ����p����"Vڦ��8�������d�]��)�;�3�|Fë�������N��ˆx���:�J\�����(hF��Ф�(Tu��qdq�@�xRw�X�h����I7���y���R�u2ؗ���ٔ��	rGT��Z�"��ܼ��(����&-]mݽ��.>N^n~��������/?O_O���/�����ܹ~��䏟�!!�Tc�pD aX��A�n�N$2bHN�|�$f�<���"��{V�"'�Y�M4���3��4��6ẖ�D�Ξ��e���1�AN]��8�-c��%���Φ�6fb�o�4r��f�h/�޽|���8���ߝ���n>�g��u�ɮ�r��,g�(Hw��J���� k�j�țeA���kd�Pw�Ӓ�샰C!k��Y�M�Z�(q�l�1�O�G��:N$M$���)��`ҡ��U�y7#�I^e3�J�o��N���X�I���tSpW�i�m��,����0�9��o�d� /GTp�i7Iw�[�f�M��,f^���b�*��b�.
�:u�ؘ5q1V#:���V��d�D?]�U�Ld2"��Q#i�DR*5�Ru�H?�4�UV�C��I����G}�\g�p��Nq�iM$nu��&�Щ����8�y|��e@�"Z���]��i�J0C��G�\6� @��SN�����$)`$ �F3O�i^�)Sڝr��\&$�/��k���
l�� jN������ [�tz�cy�Yۙ�9t��	SBVt�o�,gZ�NJ�EA����� �~�b�A����Y�fr户����x�k���-�n�?L!E"�I{_��\褝�M��vfblJm��Zyɘ҈��fI�%
㫰�G�FiY�<�@iMZ]�ǘ��ʏ8��i�۲}�e�r�\�ʙ��( LL��c�>�j���Mv�f���<Ėsc��̘��oTl[tS{X7[����[����o���y��ԗ�\:`F���s73~�m�Fx���旃R'[{~��`�#��
7c�Eƾ?!��2�(��8��	�9:Vz�9���\犼B�NUX��?}������]��E�*l}���E`\�3�~W�b>ڻ���臯B��ߏ���/����rV��~���
�?��/�T��?>���_�H�b0~�6ؕx�"۫ �@ N�~�`	OȾ:�/ ]�����;�6� 
q�D,b��r�@4X�ך87@��a��XE<�{F�"����ǋd|��XP�2vьc�W�F/��'�P��(�F<�q�߃���8
�lLc	�H>��T�Ld I�H6r�rlc	��7�`�Yx$%�XOr1[���'�x�A�/��|$#E�FC�Q��9�-�H�[�P��[	�?��2X�h*IX:r����&���^����%4�YMW�ҙ^�y�,VqR,'"X�Epv�q4����x�s��K:)b��3�J�'
�ل}
4�@�@��&q��.8��(ҁo6�Eg΂��*4�u(a�Q����-)���%�.�$��I9@�%\�ߌh'-pQJE���)J9��te��t�K_�Q ��
�)L��Γ�T�]����v�QJ��H��D�f�y���X����4�)D�zV�f���L�Bo�S�v4�j��?z���y�,�a�X��1��+��\�A���0Q`cwX�ˊ!�3a,�g=�~6���l(;�Ժ��Bafi؊��6��Šh%�A5�v�� jo(C��{���g����~����c÷��%v�ԭ�uuge%�I˻;*��aLGsϚB�*�����\�YĀR�����j��}}Q��G8���x�_�	AI��x1�*,���o����ݙjL8ȅ�ӝF�Nt�PT^7�h�6x�z>w�1l�x�0�(���|�Y�y�/���LI4�1�A���D+�ۭ02�R�g꼾���=��Hn���u���,_�L
[޼Ѷ�}7��]l�<]� ����6d�1�}8\�ҳ#�P�O�*91��i�\�����*<�ny�I�N�fe�d��u��*8Lz�j��?���p��G�۳��!1�̎���e�y��ר2����\�:m�~[w��k/�Od0~Z�e��d=�0�}ldڍ7����}��C%�8V0Ӷ}G�,iUa�Aw��(B{;�@�6T<�����BJ��iN��$�	O�հ:;�{�d�X~�}lso2LN�KQ*C��	O���bBg7y�����됋|�/��?~�_;t�Jy�!�	���
�.@Β[�!G��7`F�/���j��j|k��B*���m4��Ù���J��-uDz�n�9u�M�bݡ���Jݎȑ�r&ў%wV��13�W���}�|���'������kި���f�zܻllY��ٹ�+��7x@[�����=�X� 10��c���yj@Auf�)U}`Q`(>�8�_����;q�k���O��/�8ց�g��k;��]��}r}���o9=�<�~���f�Mp9g3�>s��X�>9���EK��X�$] �,̢qer�4LY���d�W��w�~�{k�8�Su2�v:����T����:	�u�;@�8�`�� ��`v��u(j�G(7�|�p3�'e�Fea�<�~Eh�$g}=�}��}��y.v_y�z�m�Őq��|'zz@|��p�^ hl6dr@B1�x���oHv�&�v.W�zp��yxD�9W�b[�z����c��p�k�'er�}4x��(�[�q�~��h}�h�)>�~L�t��;B�j,'w���*�~u�~����������h�Ht�a���~���}ހ�D�h�cn�f"��su�w(&�b:6x6��"x���5��ȍ�����]A������gU����`�w�U����ǅi{�����|�[���V���(����oè�9U�|c�x|�R~rs�F|Qh��(^�U(3^��|�g��6'�Kh~ݨ�+ID���u��H�r�#�S�P ����`��(|`�69tgA�n@�?�$I`��)�����9��D�|2�
w~�C'�v���?�fqW��5	Gy���	Xb!X�"R��6	h�T:Yt)9�:n)�a�ei���%�S�,<eW�g�Xr��8�v�x��wG~��,陟	=.YkU&�M8��p��cu)z�n3���h�x�6:�&`�D��s.��(v4���'}j�pG���ɜa}��
�V:�ƁO��~���(�[胭��_�q�8��i��Yr�ș臉��*�7�ۥ~<����sj�(�o�Z�Y��{Ͱ���������؋��fΈ����z����]9�J(�B���vȠ�y��I#�Y�艢)�	s�r��������X2��l�I�r�n��"&"6@a��`�y�!_�ПzUG_��pJ:p�'�����9��`9��=�@�5�ڶ]���i�:���_>�_bzlڣ�Y��_L�]�yr0��*��{��⧙�'�K	d�&9�2#ъ\fr-�
C�&�f%y'�x��]�%�P�(h-Q4]����*�����X�kvq �7�^*6�B��Qo�j����|#8��W�g��o˸�zk���**"A3m&	�
�o`b�#5C7L�A�R�%���#�*�6�w�Y�q6~����ʧ�ʮz����qgg�~���xx �GC���nI3�zx�!
�j�h��`��/�c	�A�ryTz�i2US<#zC�by��x��6�;w٩z����wi#8� ��V�����^�@�k�m(�s
�QA}�Ǥ���I�#����خO����(�rڙ��jˊ�n �z���$������%���&���&�:%R�Fb��"j<���ʪ�7&��:+�Vuc"98A��?�o;��Hi~����������*�ԊK��0'�W�A{.B�����еX�����#s�z�Q����/�5&j58�0a�P/��)s��� @�`�<�!����H�`$���!����˻`9I���X�`.6�� ?�av����in�:#�@E��gP�R�˰	�Q5�`�'���Q���Ϣ��b2P�C�1�8�P���*�L�N���ʺ���T��p�k+�"�!vi�8��@~P�W�)�v��(�������6,$���r�['���zq2:e
�yu�b��ʊ)��p)�@g�x�j6�[��#�{���=�	hi 69)!ȌQ�����'�3ۓh�My�QbǪb�n:j��1��ڷ'z�%*��&��ȉl�,�M�����d�4������������2��1!�l����ҳ�z��py-˪pʽ2�����+��7���ž0�z�V����dū�aQ�:{�3��_��1̭�j/Ss��+Ⱦ��28�N��������h����U��,!�:`;��@�{ܨ2f�S"4���_q�!�&��Rv$�{�wl��L�B,��i�'��g�jX���d�;9Zڡ�l���*���f+��76��;�t�����9�+ER� ���l�*�0��3Mӥj���x��Đ�(c�J"/6Zg�[z�*�˼�
� ��1ێ��)���S������ϝ�����UM��Ib�H��iͰ̯�I8���"�	g���@�oz��f��!)����]mʬG3����u	"}�I�Z�ɴ�P�՟��������u��J��5�����"Ҟl����*7��\�SQ�HĈ�)GR4���+�]<Q-�:���뭚x�[��ۺ]�z۝stk�s٪�-+����J�0���{
�Vرr��3P")�j�k��pܲ�ڨ�����)��4iȰ���Ǳ}�(A����򉊟7��0��N�� >�g�X'$Y�Z֓=TA�5\��BC�UZ�C��˜���B?����#��uY14A"���3�e�]�@������5Y4�\7]L��N���T�7<#E�DWuTS�䗤�Ze� 4�0XQ�IRE�
�-�TV�Z��zuEGşV$�^��cn_�Uf��=� nE�aV�U�0��Q;�R2�TRe>pN�^|��q��M�R�.T9s�RTESs]���-�)�Uc~:�>P���V?����M��E���^N�w�5U�NW�AL�<گ[�����,�'X}}nE�T��1��0JӾM�K��LɔG�~M����>J��MԞ����^J�G'��nG����I��I�NI��G���b���FmU��G�F�>��n(���w$��JH�M���ׄ�!�O͎O��+���)��I�C@8��u���k��d�@~��%���<��E!B�#B1��0��/p�`��
��=�Z��!���2/��Z:��T�^��>�����e[W��3N?.A�U�n#�*O�zZ~�9��V�UtJR���'�\���_`�iُ[�a�FZ�	���d<1����5��p�A�[mr̳�,���֘���0�O��_ˀ���'�����y���a�[��܃8��u/�(*�8B�q������<�X=+���=��϶��j�y����\�*�fЄ��G�N;M��pM���f�3<�٫6���0<��:b��D������{�a@N�Z� X��3@'�%�d�2�cy�k��s}�{��C���˜Z#TJ�6sGO C��[n׻-a'Ա�Z֘�du;�yVI��N���n�����[y�2<D\9"̻\{�L�`���伌̌�
;伳�T�#t\�X�{�3��d�K*Mk4;�>]ћ�-E���ku���->>>��c����>ڙ}!g�y*�*Zgow������7�aE?W������\
�����	e�C�F��6��X����9����	if����>&��\$�Ф� Y؄����j
-������r8AlL��CD�G�,$��'��v�f��j*g��*��X�e͞E�V�X�4�<�:N�T�Jq#8�*�_��X�&�������Ê˜�Vf ��+S�l�1�\����RdЊw�<�y�f�����I�:���Y�n�~���!1i��� �3�q4��D�V��v7�Gk��m�����]^�x��͟������>��ˣ��&�X��[�~��Q6�& ��J3���!����4�*=~VJ��Z�ɰg֫�(��AGԢ���o(�91��Nې�?�f/��!������z��B�$�H#�D���z�; _�QI��Ӱ�B�#�-�cq�b���qHs�0e�f��Qs&;��ű� �.K$5����4�c����*=i� �zr,ND�d&��4�	/m��d��i�1�:Aj�T�
E�Q���ʻ�Z}�=!���V[oŕV��Cdu5ʟs�>��:���k�"a�c�oY_��p�:0z�*h�Q-Xv�9̯�e�\H�m0�k����嬀��-` z�"V�TM!�	c8IFw�`W�3�j[�Vl�>�F�������X�]��'����\OF9e�mى^�s��;D5J�/��fhKEM1�C�Ԣ��hGN" �G]��~f��>�vco��=	�.�a;z����M��pLP��NiJmL3
,�Δ�a�����d��ET��S`�����J��5c��]�]Z�r�/������v����9b�����:��t�W�k��F��7�Fb�ڜX��BԷj�#4A��&���is�"<j�%�rw矇�Nni��*F��%�<t�3?|�Ǘ���y��{b�x�K��[���g06�Ӡ?��!IR?�T 5(I-g�JF��G��4�A��7A
��T���jѳ�ox��D8B��{�"��=N�_�Y��UAֵ�>�sV�LC�Dzӳ�d'.r�
�;@i���` h� z0��,APf��E�.:щ\�w��
�wn���'�Z�Q�P����,�Q`]�b�H%oI)��fUBBҐ';!A���8�y���5.;ثJ�:&=�I3Ћ��V�e��hȋ��-@U%V�^�d����L��J��ʦ�?�Q��C�,�b$�� ��x pm!�`��|yKP�\L�����à�nj3e��eGrBќ�7PNt��U�L�*��� @_��='�a
���� ��Y�+9=� �y���)����;���u���+`�E�	G�Egy�^#u��C�Ԥ'�I�#ȅ�L}|+ ��Ʈ��Sc�Sd���cFv��
 F�����H��A��:Ԩ�n�����%�ƋN�����������* �JS���y#\�ZG=�q�!��L��<~�Ԟ唌�J�O���X�c�.#W���u��Wǥ�W�!J5�Y��C�2��:�B�Jix�V@a�#<uHe�< [�.jrC\|�0S�o�䆨�5�TH�T��	��8�D2¦��yh�S� [�V���N/q��d&zj5�w#G�T�N�A���F@���j#�^���o����b\��ql]'�o����Fr�k�쉔s�}ig5�a���,+��(Yi�LÐV;UlVY�Q�ZV��)�鍪����Ue�rU���9L=��ڃ�I� �ɺ��
����ب�+�\̄�α�ʪ߄>�ף���E��LSLd�ao!��^�!�h7Fi6��L��vd�-�#���R����Ft����t`��0<�4�$�w��i}�P�G��0.l�*U��a�T+��J+!��UU ��K�v�ڥ%�D�ލw�Vs$�Q�zZn\2��&7�
k�w���N��{J;��]�A��u*�
��q�ց�|���	����C)d�]�9���Q����bnz�w0�����@�۶�)�+P��m���n��y�h�W|�VX>ףH�9F�C~ftR�m9$��G�^��W�"de^V����^ӊ��&���]��霑�%{��*��f�{��]�<�4�tq&D�f�b!O�k
����$(.���楼V���p:��]�{U^��h�EؓJeS���G|��+'A|����Vkצ��jm�R���R���M.�yk+���3��~~sY�&��y���Lh��Pn㻜��_�i��q7�����L�k��Dq
2�%[+�M��ܴh���+C�L��u�#Q������������j�-���Q�H�m�w�H��#>�+4
�+�C�#"�8�4��[���"�*������U!������� �.��;��9:���©�Q��:8�; �������:�����:<����H1����a|��+*��3;�A=�;������4r� j�@
��"���1�0�����7�[9� ��(���M�4"�I.~��_�W�
�"�J�=+�C�!�6�鼂C�G<?9  [`X�H�5=�5�Ђ�������aSB�a\8�e��X�]��dR=ںK�9� ����".5R�����D�8����!���>���j<��SD��;�3�|��]��V#����i6�nt7N8G>SQԻ!��``��ʔ�q��b��"�|�GC�8!��Q�6��<��&�:��!d�<���2��<5��3=�3�������$j۲�����!�B�=�J@EXA���-�:xA���搵����B��!��)3Ô��\c�uY9��H����Y���29C��T�X��\�8k�&���Er�;����=d.󻖈����/�Ǹ�K�8�c��#���˻D=������K=:=��">*/,#���\,Ǆ�=J�-���,�9,��K����8�����ȊL��L�����L���|���L�L͹R�ڌ�մ��MŜ���MȌ��ܢ�DMᬫ��M�̣�M̔����輜�4�z�zҨ�#�H��T���s�'�(턢�y-�*��J��tϰ�(��
��j�O>���|���)1��������v��D*�O��E��lυԲv�P��(m���Βxϒ� v��}b�t2r�'�T� %Oz�1B��Ot�
�(Bx��$�r�#��
����l�ћ���N R�T�r��+3�&�(�Pr�(5��'��+��%��R�Pc+���";Qv"�*�R'm'(u�&�R)�(Ux�$P	[' ��#H�!ҰT��Sa���DU�[�K�a�q��S����P%�Ԍ����.)���bIJ�TM/P�P��c�'QU�R��V���`�N�UM=����L�TuZUt��Q5�Y��]VW��%�`E�cU�ҳV�Ua��R5ַ�jM�d}�gVXuU�L�g���2Uc}�f]�h��O���@WkM�j�bM�T�VvEVrV]}�U��Xm�x��X�.�:S�r�s�s��|�TXREXW�ׄ�VnVm��~]�O�X:�S��IY��9h�I��EUٕ%�N&��T���!�Y%�P(R%M�<-v:��!Y(�ѝ����Y�И��'�	�������d=�P�K5�=�Q�:Ѥ=��G���ʆ����Lg{'u����s2Z��Psҿ$�(}':5Ya�R�uPy'�DS�ӈjϷ��v�S#�Ѽ=�8��/U\���ݧ�|��݅��T�]ܸ�Y����N\��*��������]M]���R�0����U�lN��ɤ#�DN��L؜L�ԗ|�M�$��\��m^�җ�ԣ����LN����lN�ND M����U^�MNӓ�,�D=�t�M��L�L���^�_��_�L��%���_����|��,���M��K㜫�4<ޅ�����/�8���!A��^�y�����1��c�h��EK��!���h�`��( �`>!ˡ� ��ʚ[2�(J?��j�Jܳ>!��)1�K���F��7���ԡ%�`"̊Tc�F-��C��1&cv0È��QCI�	C��*H��%D��8�h�c�����o=�N��V
�-�+D>��J�Ua��W�$h��Iz�?�(Wq3&?� U<�6J�O��Jn�v�&a��A�h�I7y
Nvc_�-<Y�DIF��T w�����Sh�\t=pBZ0�3b`�e�Sfq{ z�G^A:�4�2��o��~|��K�Yc�s�Y��!���E<Q��
^�/�)����av��#��A�&��*�-�3��~.�P&��Rֱ�.b��)
|e����bO�b��1pV�v��f~ȿ�D>�FF�ҭ��3��!8@9�v���/�eu+�n>����s? ��v��|�b���	����:�Xҟ�J�r�n8����S�=y����k�/e0�(>0*HE�G�a
�80ܝ3f�l�
	BC�0�?fZv� -��b�f�Ҋ#�#j��@��d�隣"���xI��f�FO��;k)���)�����l�ݢ�D����У��:Ӯ���������뽎�Ń��4����kc�:5h6�T�?���@�����c��@��]�-����V5�3��Fo9��We�g8�k�f1�>F�V�lj�es���b��^#(8Q�.��pW�e���jp5I����2f���g>i����%[hj�q��n;44�'c�6l�N�nf�Ķ�G�����A����F�������r����H	ʫ1��q>"�oȦ�\���젛m2��B	���r����N�/�rW���k?/�)�(t�nJ�p(�c���މW��ޥ�����?�`����"��������S�<��!&�2�@7,h�o��^��6���dK�FiQ�(w4?�Nw���MΔ�ޥ⨿�>��F�zL�5v��b��`��ڝ���pΞ�r{�)?���X�֞�?)����)�hWv��p��=��m.�
 �qc��3	}/�k,W�>w�t�$]�C�)s����`G��Cn_Wg^g���E��쎄�(�����֥\�2Q�<�6�$~����i<׃���U�xSPE�"#dS&mK�ղ�4��줗��E�6H�����C{�^M�u�$[Ҋ\�Ni �o��+�����m��3wO&;�yqI�&:DuQ�f0a��Q
�ͪT�i��J��;��bx�y��N���8'n�^�Ckqp��ğ�fO�g��d�i�r�l��Ǝ�{�*�q���s6s��|����w!�xy��hF������� μ�w"���
����'| |`��k󾿰�踨k�J�<qy���Q�s�D�9J���p�?|� �Q�����E�{Z�GO�؆�d�DH қ����̄��Y1j,f�&�/���"'� ��u��z_�	�y�ʱ�U��7ge�K��{�V ��h<M2���D��)j����-������1�l>���5�힕K�ꋾ�I�z�0}j&���� @�2��-^�$�@T2bB�0��6�8� T���V�V�q��.2�Z��
_$7�6<$�"��	��I�teZ���:�Opno���e)Aqw�Ws��k������I�"��-���[�O̦<U�!�3�a�}o.b̨q#ǎ?��hы�<c�)y�K�^=J���$��<`LE��TȠjF5�)�eb��M1,�!�ԚN��2�뉧'\�� CfQ�����t*L�歘W�("��^�0bhͻz���TcC	h�zr[!����>��}�bĎĒO�@
����T�r&�sI
������B�C���~`��ǆӱI�]��^�TE�.�	쁤y4���v;�L��2Jʉӻ�̮};��޿��3�ޞ���׹~o�VJ�J[)+�(�!�(��|G��s4c��S�Ӡ�B�`n�!1@a�D،�~ba'�t���#z
Q�(t�sQ�0tX���E��`A#^��1��%�2�h�F�8�D��!z��1^xSRY��Wb���wTW�z]v��>�	�Ul7x��\S��W,ăZPrx��8N�6M�����m�`'_u�	\	���S&�ب��v��=\ͣl(@��`�p\�-wNJ\Oȹ�_X��Ë%�lUU��Y
�Ju���j�����1J��
�/)S&��ݓ�E�bΘ���b���ێ����B�%�����_魫*u'���Z�J}x�3d���� ?��W��x)u�r�H%!A���1BX䄛�r� \<�g<!j��(�$�����'���H���q�XcR�l�s�ҜI�Q��m���*,A�[��!�K����OC���y{�I[=�~M���ĂW\{����٤%�~���P'�ؽ�=J�{��B*�{
�*�ƾ�ԝ��LC�i��ۑ��p��"���+x!e3Xf`s�l���H�6�`�JV����nGK��%��}��[�pﶜ#��i��l�f\0�����y�6��h\�%�*�Q���c���P[/��Z�PtԲ�y��n�=�;��n�o:���50��/������O � ������,L^�YW!�/�H�|��ƼQ�h�n.B`�������!��F=���1�X�˰�/��!g0tS�6������t�C���G��B°$�qA|L"���'B1�R���#Vd2=�
䬲�pEPFi�����8z3\�vd�<)�lMA� i��px\�F0�D�MMɩA����tqw~��%Y�Ab�^̕�xǂ�eL/d�A������p�3�	>+�4-:� ��Wi��',��Tgt#te(7®V��������@P�Qfj��f�(����)b3���f��X�}�I��"�F� ��x��V54������
3���.��a����}��D�?�@�rB���<��3}M3�K�=�QI-`���G��n���sd��8�,�|����lf:J y���4I٢��q	Ri��B�t��$��S�L�7��ԧBu�#ϳ����Y�o��]ٞ��R�J���`VaYS��.��	�Y�&���`�r�k-30l�pY���<@�[�4��/xշ�0ꯊ=G*Ê���18��������}�(y4�e��V�@'�.�^U��Ӣ6��E�R��*X�(����m dk���vS��H5���ޖ����oG���f
��U�p��\��V�t;T�]7��'�Q\Hp�B�n��+��Vw��mnx�)i��D��mp��X=׺(/yc�]�~�ڥ�v�ۡ�6���խ�$�_�7¦��!�_�vw���p�a���-�b{��=��^+=��6�2�����+�G��������z@j{�#w��I.�����X��N�r�5��+K��D�d��l-�SJ���\�'����j>3���dX���m�3�ߌd_,6��k�ܜ�2s��_�s���)/c��bta�g)�����=Di2�9�f3�5]�HEy�%N4�0��x��S���/dWֲ�Ŏc�!�֪4�5�{���Vd��NF���ǲV6���jX���Nv��Gmv^;�Vµ��j��۵�u�oD�n7���v�^=nmo������m�@{��^�%�|h��&Hv���y�{ଂ����I ���q���fG\��6��-�t3\����6�f�cd�8��M�oӑ��Gw�_Er�{	4'w��g��<����}>�o\�D������#�;EO7ˍm�h�j��:׻�`'������YLd⦘���ڝ��8�&�����ܴ���o_p~��>�
��',w�X�=�{o�����|?p�l�7�g0u�{��ş��G�w蒾D�?��y��ѻ��8�:�ko����:�M������޵8��xH�&�}�Yj�0��2Ug�G���/\U}��o�+̆}�4j�o�Q��A��WB��Kȿ&�]�	�(�.=�F���!Fː�����єy��^:�ޟR%-`넋0G�\euMU���d��0���p|V;``-��f� )���¿�{d��F(]ԣ\��Y��H���J�D
6�`-̊	6���^q`v�p���Rf)��đ���bH�rW� L�u�����!/) �i�������M�՜��_���0_9_�P����V�M9�� �t_&� ��sWKe�%"2���*9��U ����O��H�Z
�;�N������a-�b�M��V��N"�VyY0�W��fS��".!��`�8��T!��0c�V�� �j��<
�=
V�Rhd�'�`�Re�EfdU��| 0ي~x���4Ci�d|��F'ђ	�c3�Uq@�=:�b�@1C�8�"-��DRd�ѓ`��be��K��$�V�Y�a�dG �� �'V�!^���L���K�Q@n�#>CH�����M�"����/��AD�PQ�`ɤS��8�}�JN@��i����*��%���U�)VdZ�eԼ�#���Z*d<�UW-0N�K��'�3b��(#B�`
� B�"�N.��Y5�X� ,��k��7bH8�
Qi�ej���c���&���	T�`e��B�怦:�>j�/je4��l�cX��]&���R�a9dD*M���q"g6�e��b�͢J���[NetΐK�$��dH���}�b�Z��9��HBЋ� �'�݆ 2�߻$%'Z���Z5��{R�6�!���r�^���l(G����HX&�|��7IAR�arRh�N�r�"�'U��j��f��0zU#6^)�fn�&gڦ��Ux�x��@!�����F�iv#|�Й�&>�҈����@�cT�e#��6.�^���؟@V���� �#
V��
��p�*%��x����.Ξ���r��%Wj�\���!U��@�\��E�vV���������(�C!�F~zM�a���ġR���z:%N��{Z�T^�+��KJ�R�,�a¡ZgIv"o�"V�V�G$h��cN=�֧J�髆���i�����Rә�ޓ�j��%C��6�`<&��Nht��\)	)a�I�3���(��&'�\X-�bL�a�cٌ�'b�쀨Bv&�i���g�	U�&_��'�(�
�kfi�n���h��h��J���h�r4�
��k����r�L=h��v˜��'���*j��j���Awf�v�*)����z_�^�J�z�к6�˔P�x%!�X6�FŃ~�=����'�z���U�V���=�X���u�B�f��IdǢm�n��<d�e��&k0��?z Y��5f1r�6B�����^����I T�� �r �<���訁Z	F6tR������'�R��b��I�^t��J	��u���H�h)hb�g�ĥ��oh4e,�~��m�/���fds+��d�d� �OJ/�N��� {���^�h!��^�:�g��,a�X�:u%�v�	�Y@M�le݋>DNH�z>���[B�ԝ��rF�$�)~[��L����\ƭ�� �v��=�#��x��	���!0cd �@�&"!D/����q�F�
#H=����������'�}��)Yù��"-����.�o�m������F���.��z�L$Ҝ,��,ΰ�S�:P} 3�I�0�Xő ��4�� U�Ā��P��OT4#�M �֍$Z]�����0���h��p��%�n��n�X繒��X�f�$�n��r�����0��p��F��FK����2�b(��ȊA�2D�����dD҂�T ,y�L]����|t��4�!��:�S�٨A9"2����P�\Q�i�_���K�AAf�0E�K���ah�d��)�@�"<�P_��a�g/O��$��3�T�)@�2��r?��B����rH/�֊!(�0�� �Qe���s�O��E�c=Z��RF��guhɫm6�8N�<R'G蒠6K����2+��H/&�*)�l�5��V��<��Q2\��+e�-&pU��8�1�z�`�d��U��C�a�-C��q:tBc�F6��������I|�y�0�L�l�2�K;m�KӁ��T3�K[�#���E�[�ߌ�IXT�>mf������i�a8s-����3��Ϩ�����|�O�6��s��9)�9��vP��� �x�P��W�v�+A�.�&����*��u�%G��Mq󖉝�5�KSī}�w�lM,P��e~�c�Q�U%� s���x�#u�J�����x���h2d�t�g������_)x90�8������w�7~T�U�Ms�E�*fz.bP�B7�n�ǥuc����+�e�Jt��"�q�ԩ.�t�_k��mnW�I3���O&8��@�1����k×(�<T�'��6�In��y3X��eҌ���6��p�t�.�絚W4�8L��CѰN�<w����V�s*/����עCw�G�xE ���wJ.��Wdu9Wc"�E���R��-�ˮ�l#%T%�����K�9`McA�Ҋ�ń�`7���f�JVc<)ގ�<��r@m�����ץU��XT5�� �xU�O);���<����3
�3	�c�.�fn�Ҳg��D����;�[?'u�i�,z�S�w���^�EMO�b�9D{�xԉ_y:�LKe�3v����ְ)@N�4֬�P��&�0����I���Z䪀��FïۀJFo
�����S�R���T~2%Ӷ�nAƔ�%"��U�;��׏����F��;�'�p�5?���*J�k��Y�u2���{�[hz��8/.�P�$��0��M��<]1;7����M$��B{kI����r,5SX�:�}L�+�:1O|�#�X�j�� �K��Q`�ko�(����C�&f�v;o��mf %K!k^����.)\�~'S��ҬRtQ���;�:�b~��S,d��o��۪�uq�����W���ބE��]~����m$���݈1���������䝎('��.�������������C���V{��
>�M�/�J�ĮCrAO�V���L�?��18 +�ڎCe��[2��@4h]�Uٖ�|�a�8 ��i���v��q��^���y��������J 
��7h$+/)�� 33F=K5 BGC-KH�B,?Ycs{Ey{Kh7M1K!![E�qe>�������%���mK��m#ˁO�p�}k���{g�=���1e�i�i�E�����^2w���2���#T�0��f��%/ "�u@IJ]	��c�w��3���Q'U�2eS�U��eB�p%�8��b4�C�JGY�4%.bE��R���!��,�.{4����-z���Φ?o�ƕ;�n]�w���sHe�b`U���Y���J|O1bǍ0 �1c��,/�����εB@��Y��Ę=�N=c���2��8ٙi[���1F[��s[C��4kײC�V��i��/6�<����o;w��{v��G���v���>ϻ� ܏n�;��ɻ�F����wɯ?�l���,P	���o9О�о�󄯿�0�8$��H,��QLQ�Kt��.`�a+P�b*��q��(�,�H�� x�QG~0��`�k�\���Gx�R�l��! ; �
�L"�|4�G#��q	�`��3�3!-�o PH���$��(�t�PCG�1�/U��E�����)M��C�� 8���OAU�QI-��SQMU�UYm��Wa�U�Yi���[qU��W���׎L��_9�U3v=�Sq��4YOQ	�XT�akY��qv�h���Uf>��M�5�^@*ĭg�-[R�����
�Sr����k�ݗ�u �Yt�e��|B��׏�I�_Q���w)�؋�����f���-Ju�$���V�wv��R#�vԕ��v�i]m�c�?�`�i]fQ��9�Y{�h�?.�h����駡�Zꩩ��꫱�:eU��V�S��Z�S�xg�e	c���W"��E�_�ߥ�n��n;mq�����dnۋ�	��A�^7���UW[w�R<o��f�q 
��t'j�m;��߀D��m���ؒ9�\��s\�u/N]dNI�%[Л��t3�<����Y��{��s��7}xҝ��td��W�߇�y���r_�W�襽n���;���o����_~��N�k�eY�g�����F�p	M}����b5�.pg�X!x�eg�Z����A�-�~���7�1�,��c�*���W�����[�~E���S#s��VW��}k�.{ y����d/CZ��/riC��P�A��]��b���m��]���F���G��fFT�{m�`�:�Y���#��tW=ީL�u�W�h'G��qzBTW��w<6v/^��Q���.x�s�ć6�ɭ����o����M]�0�#�셏\�+�#�1{Dғ���fCX+q�ce-YYB�9�x����<?��tt�^S��Us��L�/1̼-1�XU�a7ӗF-����4�9љN�-�jd��̧�Z������x��q�e6K ���6x͍`}4"�
/�t��`����o�t?L�͘e�
v�t��>���YlD��X�f(�{}�n��Kw2nFtU�����)�&�LU�X����EC����Y������:�U�N���k���wՐԏ���2����i�t���+���/x��i����mS�b�?TI�r!ΘD��i�bYүʬ�1MJX΍�y]A +��JS`�z�l	�8օ�c%{�0A�җG"�����Ŵ�U{������YiJ�h3�$��V�������nI�+4��Z��8��\�.��ͥ�UM8\�ʓV_�Z5�D}R4���`L�� S�bC��#�n�G}-��z\V�a�R�j�,r�Y.�V_I�]ڄ�u'FJ	7_� >�:Ĺ��ć��Up{F��5�H�0Q<E����Ғn@��b����|*�K`���Ҧ2�k:f�1��� -ۯȾ�ܘ[҆�"Y7;���]u3�kDiY���f��߼뉨È c�gE1�1Ӥ̼�,��w#:MW$ &�ɪMfe�-ﴩ9�)yρ�� ���ʪw��+��U��Lъ4��L���,ut��|�S�dX�a�8}I�Ζy`.������:��٫$�G�iRKn�Z-.���b]�׽nߋ�x�&-�[�����eإ���]s	X�b�ȋ���1\�Fak�Gg:oֽ����H���"]3���-ߍv��d����vǲ�(��&,Q��u��و8��������!�Q�)�j���*��'t}r�����.���?k\�����MW¬C���ksmL�1�9��Ǆ����s��}�w���`���?�d��0���y7$���Զ��q�=��M^bզ��z6�?�����o]>��|��fy��w���	Cy�彿�o\V�z�Zp�N�i�:��z���k�[B���o�P���	��6�����վ[�^m�R�/[��E�c�j���6�-|��^�6�ؠ+z����7���4[���z��LT���7\p��[3ǽ��,&1O�G7b��q���ج�Ͳ5�w�����V��c�!�0�}�v�f�g����.f�ʊ*⥡�#"�bF&�6��\��(��OրK����������x�n�$k������L��\�aPj�ϧpmAΩl���	�XnS���<��g��<o���
���Ьe�TN�ԍ��-��p��������)&o�p��p�� �������.,{��&r��l�x���t���c�1������70���B�HM�A���6mnZ� �9E`4�'T�G���[rj����������
M������I���6g��<n�ZT��8��	����v��O��q��ɲG��V�� �/q[&������l&���~I�⮏01��( ��㚯�Q�1�q[��-�j�E��0��Tz1�&W�T��=%�&�!r����Y�J!Í�,��߼Ё�0�.�"�bV��F�Z:�	���R7J&W!7)��(%�+�ڭ�:"�˥��s�%��f��&'���1A1��n�_���� �eZn"�t�Uf��n�O ��,���2
�f��N�q���&o"�b�qoT�𽢯.'�mR[$�&̀0�^.�
�(������ =	�����3���#$`���
*�R1k�_�q7{�	-�����@���7k�$\��jQ����t�1/���Qs��-.��'�A��������r/�3/��*u����q��r�2=ճ��2�Ј��� �� Rk�ShR?�� S��&�S"��2��3R�P�Вd3$M��PB�p
=�[2���%ҧ��S�'�#\	�
Lc�,\D`(G��˞t�T�e�2D���!sr5�+�+��!'�9O�D��*e��N���0 ���s=��JC�=��Up������B�	3������:�4G��$�3��pN�N��N�P)v`�``d�� \��vO�:�0ۈQH3;��ԑ/1N}�5��?#�8�%��1ִ�t��KQ5U�kT�n���T�r.�>=��s5��?��[�H&���uX��X�OSt}�`�t-�ڌ0T���hROX�H�e:k/+�;��V��D��d��I���������TU�u^�U���Xp�40׊�D?BQ���'5�.S��;�&s C����8���F0)Bg�_�oOO�3y��h�:�i���OWK�aVe��L6J�T�>˯u�hd
N�o솳)	�S��@�����SS_�S3Q���d��Q%�D�"!9<��U1MuJ��5lŶ�F�U�t,�k>�TICX��e�UT�v���]̵)G�m�6IuAg����v�$-�A�c<T$3�$y�C1t��MDi���V��6C4nq��6oE�M�N�hQ�LZ�mr�5K�Vm�7�D�����rsv�[+t	��v}��V}�D�RW&]y�pk�l?��sl��y�U�����J�u1�575��S\���F*�4d[�aCo��M7�{�w/ggA��qDgeW�TѠ^�K|4�~eq�h1���2�wG=�Qo�0�)�V1��{�`A����c��8�KKQgO�P�7��'�{o6ϑLIx[%�yB8e[�{qR\�&/'sw؎�q{���qg�VC1��k�jz��y�8��z�6ؤ���fJZ.wV*v4��2�kT)�-#_�A��p?r��pq�W�w��p�JKr����X)s0{b�q�/A>L��X�֐UD��bE&.��U]Xٍ���|/>naU�-�������U�x�>9RzdP��JHYN��R��S�$%Q�d�WY�o`Mޭ�v�^�
%I�eLe�C�͘��dN��I�Dv�\�P��H�YPtٔ�9�%H�����	�����R�����8m1���Y~:��g�cr0 
�d�-B4�>��LY�BX�7n��9:��;��7#�=$�?d4 z�'��+d3H֔���8��3Z?@�d�A"�B��W:�+�飤�2T�2\�=�c;:�^zB��7*�����9x�AF��/�Al$�?���;�-�����H �"y%�U���ɺ�k��F#t
�C���:��0�bX�(ԡ"ܚ&�A����:�;����Z����B+B�
�[�;���W?a<:&�3JS꺮�̇;0���S��5O�Z-,�tNHbO�,*��#J���z(d�[|�y��躷{�)��*9��3�=y��l+�۰��+&��S{���, O�ڲ������gZՄ���͹�}���J�$���y��Oy��m��[l�A�]%录�'�K/�o9b�^`N����ky�YL ��������;�K�M�;�3 �5�I���֌�|�w��w��_G�:������5�*b��'�1�tOc|rLvc5퍡6i�`kd�T�⏅�8Xy�3�i� �T{�LȲGg��g���漊�Lk˃��<��_�-�|M��\|�<Tզz.s<�5�������˖��Vy�9����x0�ڰ���[8r��}W�Ծ������#*�[��Vx����>T���/�sG��Coq:��9}Z+��m��k@׍�j�+�����=!,�]�x����U��}کݏ�z�a�^ci��R+1z4���ű��*����s���~k�fk��k������b;s�d�ƥe���sݍE�� A3���8j$��<�����1��z����ϭ�=�J��c�D����/����W���Zz���]����ە,�ӻ�P٬X+���ӕ}$��x<��8�1�Ӌ�Yv
u���7�u���]E�*ww�nB����A��y��;��9��^��J��~�]�����׭���G7��g�������5�k�������fg�1a��o��t܀���>3u�7� �^��L�����Ǚ�:
^V���<a?_�cV�
gZ�I����^ &�~�ۅ���|��\��<~�1.����S�ݝ����I��1{?�}]������_��9C�ѯ�L��'Y�*d#�X&}�F����x�u�>����M���r_Ȳ���S}F��!@ )$��^K'�޵Y�X	6��'�qfl�ڡ����Q;ߊG�L�D������t=����4�h�����vKb�:����3YN�����~����������}kq!5D�j�weWZ��AX�KG�)T���;(�O������������74�W��'�e���(�+�Y�������������#¼���ޫ�֛����昢'K ������4���Ḙ��׆�K_�Y�r;�VM����u�W��%:o*D�Q7]���ǌ��0cʜI��͛8o�\����5��Ji##1Gﰓ�VN'��QYA����j�꿤�;mJШ\�u��c(��"�ʝ��^�`��q;
Ș(^��U�7)ZH\��!A���f�b];@�^�yv�ܺ���٧�C�M����z Q��38<]�����8u����0p�����D��qj љ��{Sǌ#t�:�c��"2����h/��Zn1e�:�$R!?�e�x��N��
0 �}�!.��삛Q#��]{�AG�8ߙb0m�[���c�`�6����I�9�N��h�(��⊗�ԙ)�(��5��ht `#B�Y[�UQM28Tc��- Y��0��(�CT�L �ep�GÄbW5$�T� P���
D� �]��%�=(�Y�y9Lai�E�Q2$�Q��dQ5�9,d!��w�0%G�qr&`_��iU.�ʒ�^V�R�� ��}����x��㗚��⭸�뮼�ǋ$���#-Y`Q�5�I��I��	�	|��	 ��
~�[(�Fc�u��^,�0Щ+�z�876�B��'?�7�;����C �0��3�}�

�����p�ﾎ�Y�R"u�0�A6\�vM��c��w��_�ީ���l5쨽���<���S�����j����z�#K��1W���V��W��¢h���4A[8u��,'�pR�\�9�əTm��V��P@w����\m�i�}e��\Xn���u���#Ψ��$�2"|T�]t�ٌ&�D��^�,�褗�+�]	���ǳX��T�2+�.��+�~�0=X��W��H�-Taw�v��,��ްe��]9f���$+t�-�����N���]��ce�/�� ��2=a�� !��%Py���x��&w��i��A�K�Tǵ���S-2�'H�
�uzj�Z�H �j��` ��'�@
W'  &dE !	[�B�P�3D!�f����__i�
r(���	)��dH�LI- 8���*��y� h@��y�EOC�������:�kW�S�(L]�cX��@�������Y�(�F�ىmw��_$)��d=㦞H�t�>��efY�h�,�GI�R����r���@��w/s�>��B�"�)(a.� 鴰y�Q���x�J��	'LaH���� �HOpơ;_s��(!(ty�h�@[_�X6�3���Cw3���� h����)0����8K�c~�sES��#> �A:���a�	;�0�"��B�`ԗ�a�=�s�6����"�3�����?��(M)�@U6��+)���0��L���A����\n��#ZO`�`�`ځkP5+�.]l@�PW�G[.�H��G8��r�C�6��+�Hɶ�B_���O��cj�2GP�A�G������@=�꒥)���հ�di�����4�*��d'{+�R�56i�|���v�"�5tY� �=�b���
*����x-O���(|$#�\^z0�̓�����%'�}���7Ӗk�+�L��A��\��k�*آ|2���e��]��8a����Q���~	�¸���f	H��g�����7]:Yni�<q8T��=�S+���
�=���'La�X�@�,ci��H�/nE4�G�m��[
W[�T���bX���GW��יB$jE+b��Dz���&&!cIi�B�*Gc0��
��\Ǌ��D`�E2��`$!P	MejK�O�"��m�jې�Z����u��B*�X&��N�f�'X�U�p{�\SX VQ���jG8�;V�.MM�'M�J��ª�� �d�^���2�oE�K�*5��z�!�v��i�ى�z����E�JM��a�	��pO�����-��KQޡz��-}����mm�^�-���9�:�k�����/�e��-�:���Gl]y�N>��H��ߌ�s��������Nf�f$�����{0��l�9�Qz6�8+ꋇ�c09�37�WŅ���`��[��;��!�P�,�RW*e���9j�ﵵ4��R��b�bm>�TڋR�ћ}�(����2Ԅ ;.%�p{�]��*�[��8��f�K�"�V��\q��C�f$��P|�ϻ����H�|�'�?��~%s��6&�1��vg�Q�8<l�;rf�<9ɍ�o�S��w2�i����K~R,��v�?{y	n\���x�qc��ޞ����	~�l{�T��K7���eNحH�0�4���/���A>.{lI��p#<�� ����+�=b���'y����3��/=x��N��7���49lYj殅V�DLTTL�rj�q�,�wB,�b&d\��L$ c#PY��wߴTäc;sDU/7�XC�4GqSrj�2v%F#G.�Ac],(T��5���qxE0�60y,�o�Yy1��I���s�d1��a�cXC�-y6a I��*WƅJ�9��h�u��A��:�fn���h�uy9v@��yy���}���|x8ؗ?v�8��|�6�����u؈�s�tx�~(��@�H���x���S��S8儉�H�����=׷�և�g����5��?0 v���R��X�kъ�ȋ�h<�Ɗ���H���芥�%�x��@�Xr�vwN�ڸ�$��Q�6g3���}'��(rR��؎tҎX�������Nq��H�(�CpB�H�$�h�� ����Ŏɐi Ɏb�&!Ac�H�	)��!!';0�Y��� �"ِ�U���\(�!9�I�x6�\�69ci4'��rRN�u�����'����h*�I਎�ғ����s�CI�	'Qu0I�%bɕ��d'9���=���YB�gi���ܓ�����W��~��Fy9 )�>鐄ٗ�x�;��YvR�ITc���iiꨓ���9c�y�;��E�%�d��ɑ�Y���y������`����������iz�ym�y��Y��y��Y�Ǜ�9�Ĺ��%�9���Nʩ���%T ��i��Ě�P��R��)�����M����ٝ��x���Y����T`՜��FoVyda�	1�i�
���y�( ���J����ש���߉��I��3 �������� �J����(Y�əp�NY�����7�*��<s��(�Ո����H.�؋8Z�6z���:J��a6���;�th��#��(��x82z��Mz-�X�>����RZ���Ȍ׷Y�&�(�}��F%^gy�@�bj��8��h|<��pJ��؇D�yX�]�8O�5�8��8�uZ84�B:�xj��p,���JJ��i���JK�rq�2*����m��}�7�j�S����_��k�$��u��U]�rU8m�Z@{��~"D��;�d�:gx1W5<4��)v2��^�<����t�B���Y5��z;X���m��Ss�ӕ,? p�c�� �m��Z��3wR�w��Rx4}fWͺ=���GtaF���dԯ�,�Z�q#*�G�gl0lO:7f�cO(H6�p>�"�R�wUuQ7W:�0L@���&��I4ζZ):�N�)����no�`#V��'���q/�h���L�3}�i�(����ko�Fy#�%� !݊��A��ą��� �~+}qQ!���S@�j�>`N�*8�@;Z��5{e~�U���
�|��1��Nl{�*n���B�REhdo\�>k}���
N��E�0+w�wִ����uJH�)zQB�(��PB(f��b��uN��>��G�vxd��WC�
�z�'�O[c�`G����mn����K�if$`&,`$a&��NC�F�{�K(QKwr�
)k��C���O��}�	�gv��*���<7�;Gfi���XX���������x�
��G��
jdk���=j=��݅Pj8���*-�*	�@woķV1��j�Rg�� ��,A���H7�f9���ɧ�O��k��\�i}<'G��
k��֩�/A8�X�e���q�#���d\�6�����LQxƻ��zgP���sZrN|a�,�)�ڶs�OАEy���JG��۷�#�^Q�����ȏ��E(x^��H!)9�W�J`;hxX���5�] �f&�#�\�M3A�Sfwllƾ�˄�#Ja�'�yɓ�%\��v]K��Ь55�-�k���
ȸZ��F�н�<΃���h��D���#/�T���8�b�����gG�� �;��֩�歙�ý��� {�C]�S��yޗJc�J<��|���j�wi�p��~l#�H?8��8(pv$E�fN���r�D�)=8�) U�PU�5h�ў��f^Rd�f:"�#@�p�eI"*ǪE�@ �[& P�O]H>@sIsfx�B=]f7�����򼾔���%UuI�D9Z`$nfI"�_�^_��LP�%�ӝ��=�v�F<�hI+fUmTH�l�Ѱ�ѡ�ђ=�W��2���Ҧ���-�����.^���Ь£k�{�
=f�º�	�g��,z���Dθ}%�
�6<�4h́�����&)�0H��Ųvd�k@�F�
x�sબ�{�}�5<o��qŏ[P����{l٬�پB����A�2��m�p.�>2^��4���N��4��#�ᲊL�{(4n��Rq74����Ω��F2��E r�a�7��izU$nK�]�����Ґ�z�A|�K�Ӊ�X��9��5��:��O[�Qk+�*Г�L�����7mB~��_����«��Dt���H�!�~� ��ڳ�R�τ@,�q�[6�Y�ɾ6��T�`|V�� ��~�g�t�������EN��Qr�#�0~?2^6�J�=>,�,�;�7J��޽�gr�#S�ߺ{S|���߁���5�-���EX�^Ž����ү�}�7l��4����!Qh��F�۰�������5�`�B�w�.q���.��^�\� N��̧-��$�,<0�o�\�K�
kb�h>	m�բ��ev.���u��V=�$	X(�Cj��o�Z�W�AvNT2g�[�G%t&�^�����Vlp���=�
-ʶ�f;���ϒp�����~�����v������
��@g�.�$��QB m�]4&��G�������f�Ƒ���Z�T��o����Ȼ�u8�DPj��D�E��^-��v�ӓ�'�ͽ�ew^�9ְ�n����������n�p���R�".�C3��C��V�$t���P�jS������w��Y����
u�2|Ǩ�߳���
��yK@Z��y�������[�Gz��~ �y��n~�-�:Q�>i{N5*݅ A�8�0T~�������	ٚ����p�T����_=���� ����/��~;����������f_�}�ީ�� 䤕����0G�4O4UW�u_��TA�l	l��u�m5c)5dR�L���v�&���f�D%�n%
����se
 ��_��G!�k	V0SJ���@�A�BA5��������Ɍ�Dʷ$C�M�N�-Q��#+<ҿ�����
I��Y��۩��""N�06_G'T8����a8Ļм�b���*����4���k�tvuˑ��y�z�{�|�}��xt����n�	_Wbch��1E6:�a�"�'bK�pcl0����䨄�f��Ec�d|t�x�NʍSX�d�g紜�V��i��*EBq����S�L�I��-�"cQ�e `��<D�,���J  bP۰�Ƿ�>�(R�@J���݃C�M�UU�I�ĕ X6;
 ��_�a��mHSB��ډr�Y3��"���*g��9��\���?	I��X�Ñꖞ�[x&i�4�ȁd��%��c���s�ѥOG�ď��d�N�����FM�� =��pڔ�����G��!��5������7T�B3�J�;q��/l�ȾXtA���� @8�<�>���P�i+`����Kl@0plb>�>������Z΋��3O@��p�?�4���A�ߋ���#����N����K0�sL2{�R��ے�'ɱ�2�nZ"\�f�/��I!%�h�nd�,%��;�'���28�j4�Ն�C�Dw�(����7%�zt��a0I���i��$@ 
�P���CM�|�SC�U�Ӫ�6R"�T,����py�T=�|,1���FB|�P�"��2O�):�&q3�Aq�k�%;��F�}4Z9�o�h$��kڌ�L�x`��^&���+�;��q��CE,.�H����bb8.v�8<.�d����UY���A���H'Q�5�S��iDHrΐ��zhB�I�V��i:hJ �Q�$`6ө�M����� ��ڙ��\BA>c~�݌ŋZ���9-���|U@�`����o�S�;K�&(o(�uqG���ϗΕtqs��mᒬ*��j�rm�ޖN�6�,#<������۾2���E;�>�&�����3�F�y��
Ȑ����!�	��Lc�mP+��<b��)�W�-�p5����JKy�}]>������.�˕�m~�8irL&8�589����D��3���^b�}�$�sͰ~>�xÊS�0��y�T���}N�8��a�\�LxB�P�4��0~�Lq-�H�$��g�	
:r�z�FA�%�<��xH.qhH��ܠ$~FM$	3m�m3G�p�"$`�gd��@a����ZF�X�(�ƥ=�i7���N�FH�g!SD�q؆�d"���d�F��@��j�0�i�m��������a���
=�IP��9�����(p(�B�d�,�JXƒB��e-mIZ�2��d+wyK`�2����*Y�Kb�ʗ�f-���g3��8�,�ٲ$,���T�4���k�2��t�0e��4�Q�$',IK	Ms �9�6eY�z6Ӛ�e;���n3����9�	N~	�&0�y�Wt��ģ1�C�R��hG=:I�M wcBW$��
ye)e�JW:��J �*��K1�R]$c Q�iW�P!��	;��Lu��H�B�,�W� 7�z%:uiS�*ԠV5�)]�CWn�՞j��`�#O�ꍘv��Z�"*ԓ�V),��R���;����h��j�ڕ�&e�UŊ��h����+�jU��u	�$��BV�|����^�U����xW��Φv�MmL�5�~U�*��P��������[Ӻ*��F���i�
�֖���͟CXKֆu�LU��.�Qx|T���nw5*��aifٌ��z������
Mڻ^��W��u�[�_�~e���}���E��/��/}��_�׿�o��`7�0�K��|�?��{ 0aڋak��a��5���7�^U�u!�W8��o��+c3��f0��b,�X�.���s+F�/=]Ld?+�.���,�gX�����o��-�W�V��Q_$�l�TF�M\f-/9��E/z˫;H�	���cw��g@��j�.I�	�F����mrg��G׹���,��Ê�Ғ��l���H���ĥ쇢�
�.V=M����Vo��`u�[Gݧ����~��!�қF֍t=o�^+U�*���^R.�V�RWܢ�IN���WP#��؞�[��>[�zut�M������v��]&�tϖ�P]k���\NC�U�n�6��@\���q�ch�2Ԗ��A.�qF\�
�6+^�Y��CWh-:q_t�(�=�Py�3n�;?�qh�3��DhCé,���ބ�C_�����B9�P�=�|��+����|���~u��M��Q�)�N%�� 9]b��	m��K�}fX�dA)i��x/�^��v�a�|E�jp��6|/r�w2Y�F%��dH��m�Dn���l�SZ�T��.��]�28㿾��Hf�t_��,%��=�@�o.z�Y�}�}���i�=�n�,z�q��\�$XuY6X�BUT�O��,�7
��QF�FE>]�҆��/~��.x9�M�W� ���Ì��D�KZ��*o4x}�ӊIR@�Q�b��Hm�>�����i�پ�8<�@�@o)��9>������+GJ�s��[�]����{�A˽��=۽��A��A{p!~Ѥ|9=b�<H���+b�J;��:�#˳�
�>���ӝ�-84�ū;`���¤Y#����%���h��㻓� ���c=2;��3�<}=���cC?1=����Y���{��Ѥ'��?a��*��=!�AL�DMD��:뚺�� �	:ń8E�H��S�ZExQ>���E����8ʢ���؄nQS!�S=)E�۔��a���(�;�B�{5��B���
̜&Y�ldF\DE_(����\1G�;�곉^�����s��������3�O��M�G��?l!K��+��{��	8<��̨	��N��)���By�\�E8J"�d?Cػ�PH�A��kȲk�qp�j�3�*|�9�F��F���J=�
=.ڢ��B�9=#��9Č���FJ��"��I)ĤO,H��J��A|�D�KJ��	L�y��VDG�K���?ST�t�!�)˰�[���i�,?b��H?\\�C ��I�ɳF���U<�w���@�zAt�\��ȁ��<���K瓞�>�K�<�������e��pl��� ��R��,L�#G�L	�E4L�\�Ge�A=�J��J��ʪN��=��A� �-��F����N<����@���N��£��$ ��e�ΐ�9D\̀��IB$B,���H�H�-̣�ʀh{�	-�I�hSC�Tr�'���NGDâLģ�I�|�a������J,N���28}�:~���KR�M��?�P�=Q����N5C_��n����d�郎	*��|LV|�4�
���7!nA�xľ������9L"P��x��c��D& ��{���!���fddA{���w)�ֳ�X�@n܆	}�3�A�	/��$�S?���=���hP�cN�|�\B+�
]CA%G��R�=.D��K�8����Ի�D��*%o9�Jd�AT¼��n1�ˋ<��@�䅋��[�Q��DUMJ�@P�T��"��H�K��G5�����4�?�VjM����AԴLMwqM��S2:�QM��DSW��V�F���,�R����>T5�a�4�ymW��S5���V^�Q�JѼ���c����t o�LZɆ�[�����!��ی�Ɍ�����cdͯ�V{)��>�LA�W�9�w�r��6�Sl�!m�V��Y�A΀PN�	E$|J(4O�����B��3Vyx˲�N��T<�$2DdK�e�C	�R,Ix [S��|C&�>Y�0��X`�UҊѵP�D��<B�lϭPd��HMB Ц���P�)��M\����D͛�Qu�Gj�l���QQ9�4%
n��9!Q��	���jŕ�%��-(I8W^iG��%v	#��ċܔ�q�ܶ��[�>�Q��%fRk�5�k�X����zٍ2�3�Au$LfzH�m��U�US�ՆٱS���u ��M_����|��%�#�T@>�\ �&"+PHZJ�E$ ���ʩ�!"6��۝(���e���9�\b`�	P�E���^�����*۩�G�\`j�8�I���m%�{�	�Z�$���%�:p�@J��8�;9�s�d������!���J=]_%^�}h\�ŗl���}��N�ׄ�D�ΌЏ�`���xщ�P��b(�l��0��E������)Æ�BvIE����U@:?��"�O�̀m�uؗ�dT�c�������ؔX��=(RL6�c�Y�96� d:�]�Y��;�>Р����\Ec[��U�����0�:��3y���Y&.fc�'�_8B)�'H$7�_i �{QH��V��(�� `@�Qp���ɫ�ۗ�֓ZդR<zPB�a�NG�߶�f�\��3�O��[��I51*b�u�6�8h *h��D4�w�Hp0; �����
����:=f�6��5�}	Qi]�yϘ�a����>T�\�8��(�m��g��� �p��Rˌ����aL~M��$F��wn��lMHN�tMM$U�W��Z�W��9�E�!_ri�u��X���	<���v���X�W�z��]	�(�V�^ڏ�k�m�#&�$.Dz��f����"rJEE�Q��8�&o��~�u���
NugL�NM�]�����ZLP�^�9V��g�}���'�dRI'�ք��g%�&��V�a�R���ƈ��!���$h�lhU��k���`�k�B��Q�$�"�^h�]��i�-n��i�i=��tEcֹ���)n�^4@��WN ��� �ec��p1�V��G^�H��X�%p���x]�T6oɉ�L�oЈe
��ٴea�Mp�Mfa�_n��\=�ki�n���d�aef�A �d��SkI���6l6����cnP�����K"8vV���T�C�%��p(�e��l�����F5��&@�V�|J
pp�|�>�*Hʴ���V�hv�Ş�9��N��>�k,oÓ�u�C;f�\o��t?�kb�k�q4��VK��|�L��U ��
��V��d��a�H��ը�S�������ߐ��=ү��`uظQ�>E�E?� ���QR Yv�R������Y�H�]H�i�m�fqsaϕ`�o�F��v�?M�ⱞ�����#BiQ�-yk7ql0ޢ��6�R�$�:��[I/xl�nG��AZ�8��%�D��S$����?J�A`�
?#���w6$��!,*��&�fA)��P`�3h<�RZt�Ϙ�@��3)M�'��"��3�RV�>�mN�v$�a��oG�x�z�B�eh�!Gh�z@�c�t|_���B�E_��7��.�6x��J'��f�.q���ca	 E.�V�_��^���D��6��)���7	gǠ"�K�0���tTjv�	�ۈYK�C����^u}dk/�L�0�شI[�#���)s8|ߡ��pj�}�@�Tٲ׿�u�ftA�g��f������{����:[�%v���3'����~�3'��S9�#�j�9i�>(����']�^���r* �g�'9�_�Y�~r�j/Κ
1�z���!�)�c˳�u$��m]��ǧ�{��n�����JR��6�p��/�����3:�^���7<.����;>�?��Y"��M`׀�� �`�b� �bd��d �%��@&�f'�g����������jh�'�+�lfG*�l�@n��-����0��(�*��n�2g�f��n������r��f��8y���3Tph�56�{:2o��6nt����p�t�
,L`5���&+�%|�<雦mݨn�a������@���#@#E&RĨ�����c�&Μ:w����'�55�T�(�I+y0�4�ʨJ���Dr��UI3Yfe�	��\��l�1��Je;��X"Z�m��(I�tc������`����:�1N{��!Õ�R�6Y���^�����̔��l������4����\Nǅ}	t`gYiK��K$�׃��PQ���Pg捕��J�k�mk:0u�z��N�oe�H���5��&U�m���߲��^���)�3=��C5 �x �	*���pl�AX!!QX ��MP���N���.�(ăX�0�\%�PĈJ�`����6l�b�f�?4Ѣ�!
�a��Dű@��C:�#�SD9�!��"�0�(2�8�ZY�$L)�� ����m��&�q�9�l��Tp�e{B�&c ����1�hPFFM}��^����h�h�)�^dZ��yJʗ��^�V�n����*)����)j}��)���ݬ�訫�����v!���	���5�l�Ĵlh���ծ�l{̶�-���,�[��(Z��+�|�{٢ ��f����b�5����멷���� $�;�}�y��ҹ0�;�0�>u�'diP�g�l0����+����/�#�wr��ƻﺏ"*l��+��+�	� ���#�\*\��z�m1�{r�CgR2�����3����^�O�������.��>[��_�l�����r�O++��2��E "��h� (�`�m42��\��8�\v�rS�e����sO��x_�Р�M���:�"�Vt�eO�8ٗ�1���Y���x�1��~;�,0�f�;�r�o�α�����r���+��:_�Ŧ~�;־ד��G�}ɓ~������%���?O20�`,���̲�u�	L���L�P9)i~���?>,0}cի�0��b�_��E0W�MS�:��6,s��q��`��;�)�uޚr'�Ұ�6����?�NO;D�*'7ieN��+�������Y����ofPbG����;]�J5��=�5;ӨF4�+i�#��օ>~�k�#�A�����3��vָ��Z�4��7�E�-�i�"��xE'��t3�[��tF��q̳��A�'z���L\X#����.��x�C>ܰ���%.i��&ϕ<�]
瀽㥡Bn�0�^K��,�u�M�/Z������:m�  �&�ՁdΛt#'�
0q��{W씝JظZua����(p�
�pa����-V
�Z�W��7�!�U[d�,�Ň^���hA�ƨ���y����������*���1c����/�ˮ岦6�)N�@E�ԇ������8J�kD]% �!ƌ�	��������R���"���eC�����Oy<+}E*���{_$��ܥ/��5�XpV�UE�5�����6�W-�%r;	�kR�,r��gC[&�$Hm#�$�" �x�.R�m��PRY	0^N�^@�Fs��ղ����EE����0P�Ci߰�4�͚`�+p�+ܳ�/Vt�7��<�� ��c�+/�Ӄ�k�[à���]^���Xt�����и����{�6����W��t�w�A5�f�[�U�8�YJ�!T���H{\���b�}0�#���.��+m�ã��Ң_h99�e�d >1���W�e�K1q��܊����$��ٹ���!Z\�Ƹ�����94ydb���	6����V��������H�`3  �)s�b�jT_0,�J^���A<sL�\�g�l�.^%�_�`�a����0�-�Q�S{��,��q���Ք�u�������sy�)i�Ϣ(��ό�k�}�.�@�EE���t|U��9�y>s1k�-��T��Z���ׁAY�^��}�V��[��k�@���7ȋn�q��lm�زm Ԛ�kT��?γ�x�n����C/Z|��tF-�y�[w�v�o�vL�r䬴X�W2��ҿ!xf'yXFq�w��`,��9^r��A0��Ir9Zವ�)�ƴ��S>q	T������V�$[���:)Ո9�\�����޷����3]b
��.c��_����:~I\ia"���	�f.�r���х�)a0����I��8<}�"I��X;��:9�}۝�r�ɾ��lD{_�$�P_���Uw���S�閿<����v���B]��AƠǜ�Z��f�
E�c;�PE��]��;9�teyM��ԧt�s�5�a��n!�cv���j��"�lTU��UF�9�+\���H��J���H6�A����\�ų׍�C����-�<��/=S^�/�ɜ.�I�~��&1iZ}�4��	�7�>Q��,`=1:y�9A;9�Jp�8�7�K�ӌ=��冬X�P�{�Q�X��\!�fS�s��ZyZU�_~����L9z6��{Q�m��XT�ɠ:�S�e���?a�b�S����<��u�~!�������}�_��qA)��MU�J_Ш���p����ܡ��!�����a���"j@^�!��_��\�X�K[��[U���$ݸXc�U�m���#zz�^�$�c������"��>���)�W�L�\���佔���с��2.��a�vq�l�����_12�T�8b)��#��tc��	~"�aGn��	�朚�%h�:�]I؊I��)�c��FW��)fc���T�T�V�d�b���7v�8��8"!]��<�X�OA� :���J#3��IH�V2��1`�ݡ8.bʤ9V�b�Y�S5
"�a�8b
* �(�����ޥ�۹'�����^I�V!�����!��Q���$���d�A�f���C6�p��a!��Q��|UB�W8�g��Q����5��_K��b.�j�d�ha�H^�Q�8@DZ�D&Z֙!���}#f�h^&hR��}�hBdŔ&h�O�i௽�2!�D�5e�=�&WEb�&>#	�O3iZ?��Q@�`���̦�%ad�#9V�&L��	� s���X
g�<Z`�G��A4�$c��{c�VO��J�$_�!��~�Z���M����QvYf7�%b�\ʥ�r�%MZf��!L�'X��%�N%�Rڞ`
:�)���c��Hmh���eY�ն=K�.>�.�d��a-%����b�cW]\��NnV,��^aF���/�_|�'�V�L)����m�}��7"����,ai�my~�7jgh�����)P�#�)������O���8j�=� ��bu�q���TF5gg��=��u�bb��6i8f��R$uvgx��zgH�	G��'nI&OA&{Z����N`)�!�N&��$Ȕ�ƥXe�=�N��nP��)��K����ѠB�Qb޹"T���9e>�ђ�[�����������%_�����-�5\�j��g~����.6߈)�]+&'����j}�a�I)�&��ڄ�����4
�~���j��[q��n,�v��r����R(~���)�\f�~����Ɗlh�&ǖ��>��z,!4��M�7�+mR�.�˾��ޗ;B*����>�9ي�r�B��&�. 
z�
"`%9 9�оl���y�@��n�n���J��b���^*̊�Ǫ,��l���-�`�����v�-�B˒���m�-�.���ml).�"��N.�V��^.�f��n.�v��~.膮�.�6lb�-��R�Z����N� �� .�nj��e�^��
@ɪm�"h�N��ڭ����~h���D���iO�) MkQmQ'%*TZ\�&��R�y��)�&�݌"�^��nX���M��̍���Ư��h]*/�����-��o�h������ˆk����&���r.G�O0W�_0�g��r��2j�>Ґ��ǽș�� I	^[����
+�Y������d]����8����0�������&M�]��071I	,1OqS��@q�p[�	�F]���>��1���1�q7�cL��K��}�G}ll[��α��)�B|Xf��۱ddkT�a�G|�n �1t�klUr$��1�� K�&�%�1=�f�~9��bt�&�$WG��b|T'�q�ib[�+/'��q�'�.#�*��r,�����~�j�z��Iز0K�2O�#�Ee��gTrw�Fgr,O-|t32o5�/��!?3Y��9�2\�.C,_sp��:c�0�D%m��ꪱ?�3@�@4A�,�$�G��%?�G<�1��3�=0CtEhDC$D���
(X�=Db�GO�o�P+@H-�F��EWVGK�Cȴ1`�D�4=l41�45��OϴP5Q?PEuO�t.�tKuE�N�BC�E,4V�q���sA5X��X�5Yo��]�g����+q[��&-1c�s9���^�\^W�r@_�`�u�I]WH)k��ր]S�_k�,��,6�X�b����pF��[�h�H���0
����kWq��j#�d��h�ph�Rq��r5�zuY�p7q7���z&.�f�W��.-�:y�,�>wǞ4p�m:�Dw�-�b�_�)�.���m���?>�uu,�' �7|����u;j|�7FZ�}�7���������{��{�}��^'����x�GxO7�|{�LE�77�o8�w��8�����8�����8�����8��q�:8?����7�C�������X��Uڸ�ʨ^no���������A�}���޻<J����x��n~N���(���Oy��k�#xW�CѶ����#y�P�86������/y�5
�3�/��	闟��sj�7���8�k8�7��?:�G��O:�W��w�AW��8�O�V78�o�u�K��C'��ۅb�y�+��4Г/�ZH7q����{�@��8z'����7tQӪ{�}��~�7��x�G�u)��dM�K�z�7�w����[��9xr�x�_:�����;�����{���O%:��;jɸ��x�b�Wx��������8�Uy��7���� b{���:YTڸ���8�h���;�Ǐ+�V�\�y��<��L�O|Uy���<Zym|�9~O@@n�V���y��s���{�o���;���=�'��/=�{�H
������v��~g�@��J����c��s9:y�����O��c{��#|ፋz��9ɓ��G���|���.�[/�?x+;�?;��7ngH�9��z�>rC��?��G���;�_>�g��o>��7�7���ꪼ��v�{��V��ȠsMz�>~�z����w֔�ٿ��?9����S�Q�|A��(M�����Ԙ߾SM��h 9_
�3?��<�۹g��$��z�	���/���竺�{}�?�ǿ�Ͽ�{�Ыz�K��������- 	´Vd��)�"�+�l�3����jR����/�]h�ߠ%2�&4ΰ���.�U��fq�.�����'ȕ�$c����f6�G�s�����ʫ����hp�m�O���12�ӑ�4Tt����5Uu�����
�)S�򲦖�"J�����w�"���X�v�Y9�ٰĸ��'��+
&jE �+E#{��F({�Y�ی����Iڹ�)�y���zQ�i�7��=����) �@�28�{��I1�ڐ̀2�Y�a�)攵��Ҡ˘���5�����{ ��屋@���0,�,\���R��UT�S�V�zkV�JFmr*+G��NA�jv�)F��,����� ^�l�K����)�@��v%����f��b�XC5s������ѣG�a����ʀ��b�E��� �m=�'�� k��up�É7~9,�c-�n�i�(�D�V'H=؉�#>��Q���/3.�p4]i����AX;Bl�	W`~���Ħ�k��ȧlI��
��?��@���n�B�[襂*�(�b�P�����eԐ���1�0q.�e���m��2&Xt��f����r�õ��䊶� ���#?�J��!�1&�y(�ܒK.���I�xOBM�\-2,����;M������p�	�B��G�l))���N�A�]��F�Q��$���d�L)���4���¨�L��K���0GD'�����/XO&�`5����Hp�V���B�4e2 �h��x�|GB C����i��WS��S��M�f�PW=v\fM�XdnV�xz�D_	�R�ɍ�H����z����
mR��$ѩ�4��:$�8M3)��b�,?��6cFrԫ�9e�Y�sA&a��h�h8.E4�E���˞��	���H9�2R>�J;.m�f$�,ZǏa���'>y裵�Z/��^Ra~�듯>��VTR��m;ɲ%0�n�0`�,��n���;��|�O�q	�.�b��{�^(ϛ����r�UU��]"����V����]) 1S��{� ���t�� Χ�x2���Ԭ�f<u�c���{�@�ׁ�of��o�������^z|>s�e����~y���o�o��v&б��wi��ޟ���GnGp�S��43�M@s�C��@Z@���]�v�>����'(�	���8x��i x)t���#��$k�ʔ�Gp0{Qs��r2��ױ :P�P�Zu�	�@D�M���"�B�AJ��9� WS��i�ٳ�@$`D�a@r���qXEF�����f&��y������	�#q��U�{z3D�	���S�HC:���Q�T5�� ��TDs%AI KJ�S�F�������B�1 ")��Iv)�\�`��Dt��d�����ѫ��˝���ݥ�C̜��<�.h�����4�1�]�wQhdO�������J�#cyL��x��Ĉ�z����م���؛����h�}��D)Zѧ��`j�h�)�ӊm���x=7!
b�� :Ң�4�P!Gx��PL�@�
y�-B��d��Aã=�im���в{�/N���b�:(V��Q�*K�j=%a����bU�V}��~�ikzU+Rq�0�"C��іQjl��^��ׂ����I� '�0����<lI�6���s��BU�8}Pz��'8!�A�X����g��OC�4@�+�5�wq�S<��_b���`~��0��=E�|豦�6e�{WȰG	Z7 ��m��t��r�N��o����c���s�˂�3_k�Ź�u`okԛX�ے�P*��`�W�����`9j�;ꌫ �(I]JS>l�	�ұ��p�(�~�U�
3�T�Em�R:�̳*ܰ�@�r8���AU_T�^� Y��̠�sYep�A�Ź�؁|��5�㖎Q�hD�st�U-2�ĭ�h��1���Yֲj���?�R�IAt��@�B/s�((��k!~(α�E�2z�6G���M3fޙ�W������n[��;��n���[vʘ�y�Aj��g��.�
��4MM�I�]��'3�.;#�ueα:j�@�W����38R���A�n������9��@��7.ԙȮ�I�e��W����Wi���A�����FP�n�^	���>��u�����l����nM��k���_�o%��6����c<D-&�8�0
n�`k��#�D�p����D�,y��ۨ[����ֈE<�7����m�m;�Ֆ��i���~+"$���X�U�z�4�b�N�͒���t5xD��<�ԥ�;�-�?�v�� �K��Z�ً�����G'��B�i�"��iR#���ȴ.}�K����7��X�}՚�^c=k�l뤪lQ�je�2�C/�$�w�2�&�u|�s���5���{�)k��:��)r6b}{̰z���z���׏��,���vt�l~���fL�����{r��Vp~ ������h���y��a�E�	�/�-��W�����ƅ|kɓ?����ө������������0 �hJ�e
� �@$S�E� �/��� ���O&�5p%0y�?�}X��L��PW�[�_cPg�� ��q��j��^p��j���ڂ��	�����ra�	
ߥ9� ր
�i��0
�I��"�P�P�pÐ���װ��A�PY@߰���I�� �P� �?����p$F�qV@�gb��%�'�+)Q/q-�3�C�;GQK�q��[���p%Z����P
oaF���
����=xqb�/	����x"}���
����Q;�q�_����p�������}q'��P�����QF`/� M��Q�Ա��d���1	� ��D
a �Qr R!#R�!+R"!�!-2#��w#?R#� ߱/�Q.R#O��%�1ב"[r���	���mR'����'�F��q쏆�/h�����}��(C�)�r�N�)� xr*�g0��%u�,�R,ǒ,�2,o)g�g�,���.�P*߯'��.�8L�ʞM�v�P���$�j��v�\&���A"M�ń��� 3�\b���|2M�N#��)@X�3���31I���E3MS5)�4m�5_S��L�Tk2a��~�@`s4;D�E	�Ba��8�3�z3� ���b8��kl��r�ðb4+�*�'- ��P�!o�I�a���aL��9��;�����0��/m����t#97����8�@Y!��3,���V�6��V��R�5E<E���rA��)A�;��t�:y�<�!��S��;R�A�4�k03tEU�\>�EM3�BG�^�.�u�E7T3�/?�G�r=�H���������8�3�S��L�p3�6D��dkN�J=�O� ���ڊt:�G>W�cp�?iL9�t��T8�O�5|���9�FtD����1W�J_(�&%܀kz���k����x �z�JGg4E;�S?uSC5P�#2gS�F5b37W��������@�FOg�V�����SV��~�EcgfNẹ��0^�"��J�5�@,I���3߀��4pI%�M�T����MmuX�4<��洿v�Vו]���Zd/C�S[�G/��RK�52!'2R�F��C]3�`K��>Ǉ3PUa�UTvaAU>VP�D�< Vb{H�TH�P�dCVEtՎ��_��9�l�uKb�9����u���=�! j@�Umxm|�d�U�"����{���dE�i�vƒ"^!*V���aSSK$�r�W06CQ�R}�P�Pe^������v�Q M���k��n�a�Vb�vT#�g6E1dR1�@�6H��p�Y�OP^�N��W�6:O��������htqI�-2�4��%r��ֳ�/sO"T�F��2 "Z@x�t�h�
9�m a�>)4��wI!e����@�q��i7�7rnH�UoKAU6D����0k�]t�k�v<� lKmOlK�m��u	�D�)o��z�~���ڗF��g��4��"
^_U�y��]��d]�\��q��A�* �+�D`�Xv=�nȜdZ�DY��v�5w�
e�Vf�yn>�S�V�4n|��)$kуb�6Tu�bZ��[%x4(Xzs�;X3v+��7����W~��W�X1U�U�lja�pX��Io�q��ʀn���z��T΂��'��J�T��.N��H1\�f!�n=����ĘXgK�%��f�?���+�h�>x�,����h���q����,�n�*0��I�Um����x�j�mH�[9@a�y=�zN�L������f`]�)s��;����*�/g�KH��n��R���(<t��R`)�����yό���+� �剖�y��양��YS4+��ٔ#/��9�"w�aS�������e��>�W]]���2�*�Iw�!��-���x����He�@���-��� ��L���ܘ�/:jKz�=:q\O��itl��X��HF�(��X���C��^z��8��3IEY��N�J9�G��B(�
98���Z���UA�p96�"O��y��L�4	{��=�X�y�����~AqHK��rr�w�͇u��
ʬŹ̌��к�Iի��}9�)����Y͜�)������e	[���ՠ˯���C��Xi��xz�C�[���w�YL����z��Y{�*��Q��T��W�5̓�sE
`�O7�C�%�uO��f�-�[�4�u���d6���; �{�G�y�EY�rZ�S{�Vۧ}̧�3�m���ݬ�aZ�e��(Τ� �:��o��U��qE��Տy��c�e��;����ɉ�s9��yB⺷���#�S1�𜮭wXι�۩�Q�\��:��lp|�ə�k�z�+���ŝ�y�W<�Yܞ��w��o(��0����Xi_�@=���|�x�SJ��ӥU۽�{����e�Z��!:qUZ�w;��{�*��홃g���$��{�ߛ˿��ټ��������L����w������،}�al{��[I�����q����������W�Ȭ�e�n���bɲ/n�x�CMeӝY�'�[ȝY�Qs�$�~<z�<�ex^��%��ܱ��L�{��L�-����ؙB���s��=��؄V}�_������,��r8[p�����d�ە�+RمO�X]���}�wL���HZ�M��W��������ϼ��<:ê�����ۨɜf��r��!����=�a;/���>ݿm�g�~�'^�����=�՛�)����iZ��.���]ۚ�ž�������˷-s^�w��{���^臞���{�5�
��c��	��=f^�pjR&E��C�'�&�%�n�o��?� ��������_2$c���Y7R˞��$��#y���q$#��'R�) s���7��5��������������Þ!I�]�>"%?�y�>%���%�5���~�Q����{џ����e��^o��!����_����������_����������_����������_��������_�W������8�}�k_���Y~����_����������_����]�
���Z�޼���H�扦�ʶ�w�*L�tw���o�ņĢ�L*�̦�	�J��*��e?>�V'4ͬ���N�Gc�Ϋ����lx�������(���E7tG�6��)��h�eB��8��	*:JZzY�*�Y���Ri:K[k�!K������u+<L\l|����i�ɬ���<M]%-�����l.>N^�]�����m�����*������W>.����0�Bq�6�+hp��ĉ+Z��0�C`�]���7W��2�ʕ,5��Ub
�-kڴq#;u7{��	�VNg;==�TI!��L
5�ԩS����4"խ\)��h�dV�]˚=�6�X0��>M�&M�$�Ɍ�7�ީ/1���v���s9岶��Ō[<�����+�+��*G�0-{����{������b�QN;��>�3!���ټE��}��������w���̍A�8w��ԫ�xn8�i��O)o
�l����_������v_���50����ۯ��m����qo�q���������R`+�}^��O�e�]�2�y�������c�T�v)�(A�z#3&c��������2��"A��d�,�d�N>	e�RNIe�V^�e�Zn�e�^~	f�b�If�f��f�j��f�n�	�IΙ$�k��C�(^+t0��0�
h���h��>�h��N�(��Z*i��^�i��~�i����)���*j����j����j����*���*k��޺k�����k���+��+l������
�d0��yr��h'�f� �~{��6;.��&{n�讫n�供.����n���{o���o����/����-ݒ����^[]�Fvh��o��+p�_�q��1���q�&�,r�(��r��N��5ڣ0�'f��s�J�:��r�,�r�@���D�t�L?�t�NK�r�`��drwd��_M���1GqPO�v�j��6�l��v�i�=��m׍��0�-6�4�5��ٟ˼�7�w/��x�v;���GN9�[^�����f�3ׁc�0�����˨@�y묿~9��N�춻^;�w�y�`�ܣK`W;:�_���W� ���7}���.}��_����[���W�r�?88F�����O�=�쿿~����~���l|��y��x���t�K��E���/����@J�����$p ���b8��`�� 	+x��p�%l!
A�:�w�q;x-u�p�랷X�B�P�@b�h�$QQ�C\���t��ptr	���>"j�Kܢ��E.�q���"��7#��l�T\Q�
�3�!��_���0摎z��6��C4i�l\�*�:�)N�l�#	�HJr����%/��Ljr�KR�"�b�BvgE�)O�m�9*_(Y	�X.䃲l��W�\��:\�w� Zs�ĜFQL��l�3M�J9H�:&5���@S|��O4?��p�S�'y�7s�s�d�&;�CJB�s��T��ٰ[����g��O�0|-�A���54.�T�B
Q	��xEK<Zь������4W��$�'@�YR��̓J�K_
Ә�t�4��Mo�Ӝ���s�eJ��R��Zw�cQ��ԣ*u�K5*SS�?�P�?�
� 	��>թ\�jW��հ�u��"����QTu*���G�խ�U�d��]�z׺^qc�+��֤լ>��a�zX�*V��Mlc%�D�]0x�,T��V�f�u�g�Ά�����JU��h$_?+�ؖv����lk�T��q��U�OK�$ե��-�m�k����{�]��X������*r����j����.v�f5�f���]Lֆ������]o{�����+���y�+�:��`�X�����{`���,u���<�CX��������7��K�X�Gx����I,bF����`���-�4>q�Ql��q�e�]����W�9.�o�d'��*Kp{
���:������,ky�\1��G��c.��qq�4�y�)�(���8���r������:�y�|=��?zЄ6B���D+���n��=�CCz�A�4�a�Kk�f��F�;� �:����S�S�� � �U�ѥ:�V @�$`kZ�ZG�޵^��W�z�(�5��`�`{�26���l ��������}�hO��6ϵ�=�V���V�!A W�{���6�Y��m�{޳q7�;�jy�:���wl����:�/x���#|/8�����Y�S�����A��8�)��	x|�y�EN�<�+Oy�ctr������y�gns��\�9�9�Q�s���-�9с>t�}�G�ѕ���}�.o�͓>��3�N�zֻ^u�_]�W�zʭ��]�a��ؽ�v��]�i�x�}�����t�{�������q{�O�K�ᯆx���4��Ҏ��/?�W`ܘ��?�Ћ~��/��O��ԫ~��o��_���~�����o����~��������/����+��o����K�ԯ������k����������/��Ϗ���E��o���������������������(�H�h���	��Ȁ��(�H�h��a  ;