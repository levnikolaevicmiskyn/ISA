

package simconsts is
	constant NPIPE : integer := 4;
	constant FIXED_PIPE: integer := 5;
end simconsts;

package body simconsts is
end simconsts;
