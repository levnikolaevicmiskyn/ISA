library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MBE is
	generic(N:integer := 32);
	port(
		m_and, m_ier: in std_logic_vector(N-1 downto 0);
		z: out std_logic_vector(2*N-1 downto 0)
		);
end entity MBE;

architecture RTL of MBE is

component FA is
port(a, b, cin: in std_logic;
	s, cout: out std_logic);
end component;

component HA is
port(a, b: in std_logic;
	s, cout: out std_logic);
end component;
type matype is array(N/2 downto 0) of std_logic_vector(N downto 0); -- N/2 operands
signal pprod: matype;
signal a, a2, a_neg, a2_neg: std_logic_vector(N downto 0);
signal S: std_logic_vector(N/2 downto 0);
signal res_a, res_b: std_logic_vector(2*N-1 downto 0); 
 
-- BEGIN AUTOGEN DECL
signal st1col1: std_logic_vector(2-1 downto 0);
signal st1col2: std_logic_vector(1-1 downto 0);
signal st1col3: std_logic_vector(2-1 downto 0);
signal st1col4: std_logic_vector(2-1 downto 0);
signal st1col5: std_logic_vector(2-1 downto 0);
signal st1col6: std_logic_vector(2-1 downto 0);
signal st1col7: std_logic_vector(2-1 downto 0);
signal st1col8: std_logic_vector(2-1 downto 0);
signal st1col9: std_logic_vector(2-1 downto 0);
signal st1col10: std_logic_vector(2-1 downto 0);
signal st1col11: std_logic_vector(2-1 downto 0);
signal st1col12: std_logic_vector(2-1 downto 0);
signal st1col13: std_logic_vector(2-1 downto 0);
signal st1col14: std_logic_vector(2-1 downto 0);
signal st1col15: std_logic_vector(2-1 downto 0);
signal st1col16: std_logic_vector(2-1 downto 0);
signal st1col17: std_logic_vector(2-1 downto 0);
signal st1col18: std_logic_vector(2-1 downto 0);
signal st1col19: std_logic_vector(2-1 downto 0);
signal st1col20: std_logic_vector(2-1 downto 0);
signal st1col21: std_logic_vector(2-1 downto 0);
signal st1col22: std_logic_vector(2-1 downto 0);
signal st1col23: std_logic_vector(2-1 downto 0);
signal st1col24: std_logic_vector(2-1 downto 0);
signal st1col25: std_logic_vector(2-1 downto 0);
signal st1col26: std_logic_vector(2-1 downto 0);
signal st1col27: std_logic_vector(2-1 downto 0);
signal st1col28: std_logic_vector(2-1 downto 0);
signal st1col29: std_logic_vector(2-1 downto 0);
signal st1col30: std_logic_vector(2-1 downto 0);
signal st1col31: std_logic_vector(2-1 downto 0);
signal st1col32: std_logic_vector(2-1 downto 0);
signal st1col33: std_logic_vector(2-1 downto 0);
signal st1col34: std_logic_vector(2-1 downto 0);
signal st1col35: std_logic_vector(2-1 downto 0);
signal st1col36: std_logic_vector(2-1 downto 0);
signal st1col37: std_logic_vector(2-1 downto 0);
signal st1col38: std_logic_vector(2-1 downto 0);
signal st1col39: std_logic_vector(2-1 downto 0);
signal st1col40: std_logic_vector(2-1 downto 0);
signal st1col41: std_logic_vector(2-1 downto 0);
signal st1col42: std_logic_vector(2-1 downto 0);
signal st1col43: std_logic_vector(2-1 downto 0);
signal st1col44: std_logic_vector(2-1 downto 0);
signal st1col45: std_logic_vector(2-1 downto 0);
signal st1col46: std_logic_vector(2-1 downto 0);
signal st1col47: std_logic_vector(2-1 downto 0);
signal st1col48: std_logic_vector(2-1 downto 0);
signal st1col49: std_logic_vector(2-1 downto 0);
signal st1col50: std_logic_vector(2-1 downto 0);
signal st1col51: std_logic_vector(2-1 downto 0);
signal st1col52: std_logic_vector(2-1 downto 0);
signal st1col53: std_logic_vector(2-1 downto 0);
signal st1col54: std_logic_vector(2-1 downto 0);
signal st1col55: std_logic_vector(2-1 downto 0);
signal st1col56: std_logic_vector(2-1 downto 0);
signal st1col57: std_logic_vector(2-1 downto 0);
signal st1col58: std_logic_vector(2-1 downto 0);
signal st1col59: std_logic_vector(2-1 downto 0);
signal st1col60: std_logic_vector(2-1 downto 0);
signal st1col61: std_logic_vector(2-1 downto 0);
signal st1col62: std_logic_vector(2-1 downto 0);
signal st1col63: std_logic_vector(2-1 downto 0);
signal st1col64: std_logic_vector(2-1 downto 0);
signal st2col1: std_logic_vector(2-1 downto 0);
signal st2col2: std_logic_vector(1-1 downto 0);
signal st2col3: std_logic_vector(3-1 downto 0);
signal st2col4: std_logic_vector(2-1 downto 0);
signal st2col5: std_logic_vector(3-1 downto 0);
signal st2col6: std_logic_vector(3-1 downto 0);
signal st2col7: std_logic_vector(3-1 downto 0);
signal st2col8: std_logic_vector(3-1 downto 0);
signal st2col9: std_logic_vector(3-1 downto 0);
signal st2col10: std_logic_vector(3-1 downto 0);
signal st2col11: std_logic_vector(3-1 downto 0);
signal st2col12: std_logic_vector(3-1 downto 0);
signal st2col13: std_logic_vector(3-1 downto 0);
signal st2col14: std_logic_vector(3-1 downto 0);
signal st2col15: std_logic_vector(3-1 downto 0);
signal st2col16: std_logic_vector(3-1 downto 0);
signal st2col17: std_logic_vector(3-1 downto 0);
signal st2col18: std_logic_vector(3-1 downto 0);
signal st2col19: std_logic_vector(3-1 downto 0);
signal st2col20: std_logic_vector(3-1 downto 0);
signal st2col21: std_logic_vector(3-1 downto 0);
signal st2col22: std_logic_vector(3-1 downto 0);
signal st2col23: std_logic_vector(3-1 downto 0);
signal st2col24: std_logic_vector(3-1 downto 0);
signal st2col25: std_logic_vector(3-1 downto 0);
signal st2col26: std_logic_vector(3-1 downto 0);
signal st2col27: std_logic_vector(3-1 downto 0);
signal st2col28: std_logic_vector(3-1 downto 0);
signal st2col29: std_logic_vector(3-1 downto 0);
signal st2col30: std_logic_vector(3-1 downto 0);
signal st2col31: std_logic_vector(3-1 downto 0);
signal st2col32: std_logic_vector(3-1 downto 0);
signal st2col33: std_logic_vector(3-1 downto 0);
signal st2col34: std_logic_vector(3-1 downto 0);
signal st2col35: std_logic_vector(3-1 downto 0);
signal st2col36: std_logic_vector(3-1 downto 0);
signal st2col37: std_logic_vector(3-1 downto 0);
signal st2col38: std_logic_vector(3-1 downto 0);
signal st2col39: std_logic_vector(3-1 downto 0);
signal st2col40: std_logic_vector(3-1 downto 0);
signal st2col41: std_logic_vector(3-1 downto 0);
signal st2col42: std_logic_vector(3-1 downto 0);
signal st2col43: std_logic_vector(3-1 downto 0);
signal st2col44: std_logic_vector(3-1 downto 0);
signal st2col45: std_logic_vector(3-1 downto 0);
signal st2col46: std_logic_vector(3-1 downto 0);
signal st2col47: std_logic_vector(3-1 downto 0);
signal st2col48: std_logic_vector(3-1 downto 0);
signal st2col49: std_logic_vector(3-1 downto 0);
signal st2col50: std_logic_vector(3-1 downto 0);
signal st2col51: std_logic_vector(3-1 downto 0);
signal st2col52: std_logic_vector(3-1 downto 0);
signal st2col53: std_logic_vector(3-1 downto 0);
signal st2col54: std_logic_vector(3-1 downto 0);
signal st2col55: std_logic_vector(3-1 downto 0);
signal st2col56: std_logic_vector(3-1 downto 0);
signal st2col57: std_logic_vector(3-1 downto 0);
signal st2col58: std_logic_vector(3-1 downto 0);
signal st2col59: std_logic_vector(3-1 downto 0);
signal st2col60: std_logic_vector(3-1 downto 0);
signal st2col61: std_logic_vector(3-1 downto 0);
signal st2col62: std_logic_vector(3-1 downto 0);
signal st2col63: std_logic_vector(3-1 downto 0);
signal st2col64: std_logic_vector(3-1 downto 0);
signal st3col1: std_logic_vector(2-1 downto 0);
signal st3col2: std_logic_vector(1-1 downto 0);
signal st3col3: std_logic_vector(3-1 downto 0);
signal st3col4: std_logic_vector(2-1 downto 0);
signal st3col5: std_logic_vector(4-1 downto 0);
signal st3col6: std_logic_vector(3-1 downto 0);
signal st3col7: std_logic_vector(4-1 downto 0);
signal st3col8: std_logic_vector(4-1 downto 0);
signal st3col9: std_logic_vector(4-1 downto 0);
signal st3col10: std_logic_vector(4-1 downto 0);
signal st3col11: std_logic_vector(4-1 downto 0);
signal st3col12: std_logic_vector(4-1 downto 0);
signal st3col13: std_logic_vector(4-1 downto 0);
signal st3col14: std_logic_vector(4-1 downto 0);
signal st3col15: std_logic_vector(4-1 downto 0);
signal st3col16: std_logic_vector(4-1 downto 0);
signal st3col17: std_logic_vector(4-1 downto 0);
signal st3col18: std_logic_vector(4-1 downto 0);
signal st3col19: std_logic_vector(4-1 downto 0);
signal st3col20: std_logic_vector(4-1 downto 0);
signal st3col21: std_logic_vector(4-1 downto 0);
signal st3col22: std_logic_vector(4-1 downto 0);
signal st3col23: std_logic_vector(4-1 downto 0);
signal st3col24: std_logic_vector(4-1 downto 0);
signal st3col25: std_logic_vector(4-1 downto 0);
signal st3col26: std_logic_vector(4-1 downto 0);
signal st3col27: std_logic_vector(4-1 downto 0);
signal st3col28: std_logic_vector(4-1 downto 0);
signal st3col29: std_logic_vector(4-1 downto 0);
signal st3col30: std_logic_vector(4-1 downto 0);
signal st3col31: std_logic_vector(4-1 downto 0);
signal st3col32: std_logic_vector(4-1 downto 0);
signal st3col33: std_logic_vector(4-1 downto 0);
signal st3col34: std_logic_vector(4-1 downto 0);
signal st3col35: std_logic_vector(4-1 downto 0);
signal st3col36: std_logic_vector(4-1 downto 0);
signal st3col37: std_logic_vector(4-1 downto 0);
signal st3col38: std_logic_vector(4-1 downto 0);
signal st3col39: std_logic_vector(4-1 downto 0);
signal st3col40: std_logic_vector(4-1 downto 0);
signal st3col41: std_logic_vector(4-1 downto 0);
signal st3col42: std_logic_vector(4-1 downto 0);
signal st3col43: std_logic_vector(4-1 downto 0);
signal st3col44: std_logic_vector(4-1 downto 0);
signal st3col45: std_logic_vector(4-1 downto 0);
signal st3col46: std_logic_vector(4-1 downto 0);
signal st3col47: std_logic_vector(4-1 downto 0);
signal st3col48: std_logic_vector(4-1 downto 0);
signal st3col49: std_logic_vector(4-1 downto 0);
signal st3col50: std_logic_vector(4-1 downto 0);
signal st3col51: std_logic_vector(4-1 downto 0);
signal st3col52: std_logic_vector(4-1 downto 0);
signal st3col53: std_logic_vector(4-1 downto 0);
signal st3col54: std_logic_vector(4-1 downto 0);
signal st3col55: std_logic_vector(4-1 downto 0);
signal st3col56: std_logic_vector(4-1 downto 0);
signal st3col57: std_logic_vector(4-1 downto 0);
signal st3col58: std_logic_vector(4-1 downto 0);
signal st3col59: std_logic_vector(4-1 downto 0);
signal st3col60: std_logic_vector(4-1 downto 0);
signal st3col61: std_logic_vector(4-1 downto 0);
signal st3col62: std_logic_vector(4-1 downto 0);
signal st3col63: std_logic_vector(3-1 downto 0);
signal st3col64: std_logic_vector(2-1 downto 0);
signal st4col1: std_logic_vector(2-1 downto 0);
signal st4col2: std_logic_vector(1-1 downto 0);
signal st4col3: std_logic_vector(3-1 downto 0);
signal st4col4: std_logic_vector(2-1 downto 0);
signal st4col5: std_logic_vector(4-1 downto 0);
signal st4col6: std_logic_vector(3-1 downto 0);
signal st4col7: std_logic_vector(5-1 downto 0);
signal st4col8: std_logic_vector(4-1 downto 0);
signal st4col9: std_logic_vector(6-1 downto 0);
signal st4col10: std_logic_vector(5-1 downto 0);
signal st4col11: std_logic_vector(6-1 downto 0);
signal st4col12: std_logic_vector(6-1 downto 0);
signal st4col13: std_logic_vector(6-1 downto 0);
signal st4col14: std_logic_vector(6-1 downto 0);
signal st4col15: std_logic_vector(6-1 downto 0);
signal st4col16: std_logic_vector(6-1 downto 0);
signal st4col17: std_logic_vector(6-1 downto 0);
signal st4col18: std_logic_vector(6-1 downto 0);
signal st4col19: std_logic_vector(6-1 downto 0);
signal st4col20: std_logic_vector(6-1 downto 0);
signal st4col21: std_logic_vector(6-1 downto 0);
signal st4col22: std_logic_vector(6-1 downto 0);
signal st4col23: std_logic_vector(6-1 downto 0);
signal st4col24: std_logic_vector(6-1 downto 0);
signal st4col25: std_logic_vector(6-1 downto 0);
signal st4col26: std_logic_vector(6-1 downto 0);
signal st4col27: std_logic_vector(6-1 downto 0);
signal st4col28: std_logic_vector(6-1 downto 0);
signal st4col29: std_logic_vector(6-1 downto 0);
signal st4col30: std_logic_vector(6-1 downto 0);
signal st4col31: std_logic_vector(6-1 downto 0);
signal st4col32: std_logic_vector(6-1 downto 0);
signal st4col33: std_logic_vector(6-1 downto 0);
signal st4col34: std_logic_vector(6-1 downto 0);
signal st4col35: std_logic_vector(6-1 downto 0);
signal st4col36: std_logic_vector(6-1 downto 0);
signal st4col37: std_logic_vector(6-1 downto 0);
signal st4col38: std_logic_vector(6-1 downto 0);
signal st4col39: std_logic_vector(6-1 downto 0);
signal st4col40: std_logic_vector(6-1 downto 0);
signal st4col41: std_logic_vector(6-1 downto 0);
signal st4col42: std_logic_vector(6-1 downto 0);
signal st4col43: std_logic_vector(6-1 downto 0);
signal st4col44: std_logic_vector(6-1 downto 0);
signal st4col45: std_logic_vector(6-1 downto 0);
signal st4col46: std_logic_vector(6-1 downto 0);
signal st4col47: std_logic_vector(6-1 downto 0);
signal st4col48: std_logic_vector(6-1 downto 0);
signal st4col49: std_logic_vector(6-1 downto 0);
signal st4col50: std_logic_vector(6-1 downto 0);
signal st4col51: std_logic_vector(6-1 downto 0);
signal st4col52: std_logic_vector(6-1 downto 0);
signal st4col53: std_logic_vector(6-1 downto 0);
signal st4col54: std_logic_vector(6-1 downto 0);
signal st4col55: std_logic_vector(6-1 downto 0);
signal st4col56: std_logic_vector(6-1 downto 0);
signal st4col57: std_logic_vector(6-1 downto 0);
signal st4col58: std_logic_vector(6-1 downto 0);
signal st4col59: std_logic_vector(5-1 downto 0);
signal st4col60: std_logic_vector(4-1 downto 0);
signal st4col61: std_logic_vector(4-1 downto 0);
signal st4col62: std_logic_vector(3-1 downto 0);
signal st4col63: std_logic_vector(3-1 downto 0);
signal st4col64: std_logic_vector(2-1 downto 0);
signal st5col1: std_logic_vector(2-1 downto 0);
signal st5col2: std_logic_vector(1-1 downto 0);
signal st5col3: std_logic_vector(3-1 downto 0);
signal st5col4: std_logic_vector(2-1 downto 0);
signal st5col5: std_logic_vector(4-1 downto 0);
signal st5col6: std_logic_vector(3-1 downto 0);
signal st5col7: std_logic_vector(5-1 downto 0);
signal st5col8: std_logic_vector(4-1 downto 0);
signal st5col9: std_logic_vector(6-1 downto 0);
signal st5col10: std_logic_vector(5-1 downto 0);
signal st5col11: std_logic_vector(7-1 downto 0);
signal st5col12: std_logic_vector(6-1 downto 0);
signal st5col13: std_logic_vector(8-1 downto 0);
signal st5col14: std_logic_vector(7-1 downto 0);
signal st5col15: std_logic_vector(9-1 downto 0);
signal st5col16: std_logic_vector(8-1 downto 0);
signal st5col17: std_logic_vector(9-1 downto 0);
signal st5col18: std_logic_vector(9-1 downto 0);
signal st5col19: std_logic_vector(9-1 downto 0);
signal st5col20: std_logic_vector(9-1 downto 0);
signal st5col21: std_logic_vector(9-1 downto 0);
signal st5col22: std_logic_vector(9-1 downto 0);
signal st5col23: std_logic_vector(9-1 downto 0);
signal st5col24: std_logic_vector(9-1 downto 0);
signal st5col25: std_logic_vector(9-1 downto 0);
signal st5col26: std_logic_vector(9-1 downto 0);
signal st5col27: std_logic_vector(9-1 downto 0);
signal st5col28: std_logic_vector(9-1 downto 0);
signal st5col29: std_logic_vector(9-1 downto 0);
signal st5col30: std_logic_vector(9-1 downto 0);
signal st5col31: std_logic_vector(9-1 downto 0);
signal st5col32: std_logic_vector(9-1 downto 0);
signal st5col33: std_logic_vector(9-1 downto 0);
signal st5col34: std_logic_vector(9-1 downto 0);
signal st5col35: std_logic_vector(9-1 downto 0);
signal st5col36: std_logic_vector(9-1 downto 0);
signal st5col37: std_logic_vector(9-1 downto 0);
signal st5col38: std_logic_vector(9-1 downto 0);
signal st5col39: std_logic_vector(9-1 downto 0);
signal st5col40: std_logic_vector(9-1 downto 0);
signal st5col41: std_logic_vector(9-1 downto 0);
signal st5col42: std_logic_vector(9-1 downto 0);
signal st5col43: std_logic_vector(9-1 downto 0);
signal st5col44: std_logic_vector(9-1 downto 0);
signal st5col45: std_logic_vector(9-1 downto 0);
signal st5col46: std_logic_vector(9-1 downto 0);
signal st5col47: std_logic_vector(9-1 downto 0);
signal st5col48: std_logic_vector(9-1 downto 0);
signal st5col49: std_logic_vector(9-1 downto 0);
signal st5col50: std_logic_vector(9-1 downto 0);
signal st5col51: std_logic_vector(9-1 downto 0);
signal st5col52: std_logic_vector(9-1 downto 0);
signal st5col53: std_logic_vector(8-1 downto 0);
signal st5col54: std_logic_vector(7-1 downto 0);
signal st5col55: std_logic_vector(7-1 downto 0);
signal st5col56: std_logic_vector(6-1 downto 0);
signal st5col57: std_logic_vector(6-1 downto 0);
signal st5col58: std_logic_vector(5-1 downto 0);
signal st5col59: std_logic_vector(5-1 downto 0);
signal st5col60: std_logic_vector(4-1 downto 0);
signal st5col61: std_logic_vector(4-1 downto 0);
signal st5col62: std_logic_vector(3-1 downto 0);
signal st5col63: std_logic_vector(3-1 downto 0);
signal st5col64: std_logic_vector(2-1 downto 0);
signal st6col1: std_logic_vector(2-1 downto 0);
signal st6col2: std_logic_vector(1-1 downto 0);
signal st6col3: std_logic_vector(3-1 downto 0);
signal st6col4: std_logic_vector(2-1 downto 0);
signal st6col5: std_logic_vector(4-1 downto 0);
signal st6col6: std_logic_vector(3-1 downto 0);
signal st6col7: std_logic_vector(5-1 downto 0);
signal st6col8: std_logic_vector(4-1 downto 0);
signal st6col9: std_logic_vector(6-1 downto 0);
signal st6col10: std_logic_vector(5-1 downto 0);
signal st6col11: std_logic_vector(7-1 downto 0);
signal st6col12: std_logic_vector(6-1 downto 0);
signal st6col13: std_logic_vector(8-1 downto 0);
signal st6col14: std_logic_vector(7-1 downto 0);
signal st6col15: std_logic_vector(9-1 downto 0);
signal st6col16: std_logic_vector(8-1 downto 0);
signal st6col17: std_logic_vector(10-1 downto 0);
signal st6col18: std_logic_vector(9-1 downto 0);
signal st6col19: std_logic_vector(11-1 downto 0);
signal st6col20: std_logic_vector(10-1 downto 0);
signal st6col21: std_logic_vector(12-1 downto 0);
signal st6col22: std_logic_vector(11-1 downto 0);
signal st6col23: std_logic_vector(13-1 downto 0);
signal st6col24: std_logic_vector(12-1 downto 0);
signal st6col25: std_logic_vector(13-1 downto 0);
signal st6col26: std_logic_vector(13-1 downto 0);
signal st6col27: std_logic_vector(13-1 downto 0);
signal st6col28: std_logic_vector(13-1 downto 0);
signal st6col29: std_logic_vector(13-1 downto 0);
signal st6col30: std_logic_vector(13-1 downto 0);
signal st6col31: std_logic_vector(13-1 downto 0);
signal st6col32: std_logic_vector(13-1 downto 0);
signal st6col33: std_logic_vector(13-1 downto 0);
signal st6col34: std_logic_vector(13-1 downto 0);
signal st6col35: std_logic_vector(13-1 downto 0);
signal st6col36: std_logic_vector(13-1 downto 0);
signal st6col37: std_logic_vector(13-1 downto 0);
signal st6col38: std_logic_vector(13-1 downto 0);
signal st6col39: std_logic_vector(13-1 downto 0);
signal st6col40: std_logic_vector(13-1 downto 0);
signal st6col41: std_logic_vector(13-1 downto 0);
signal st6col42: std_logic_vector(13-1 downto 0);
signal st6col43: std_logic_vector(13-1 downto 0);
signal st6col44: std_logic_vector(13-1 downto 0);
signal st6col45: std_logic_vector(12-1 downto 0);
signal st6col46: std_logic_vector(11-1 downto 0);
signal st6col47: std_logic_vector(11-1 downto 0);
signal st6col48: std_logic_vector(10-1 downto 0);
signal st6col49: std_logic_vector(10-1 downto 0);
signal st6col50: std_logic_vector(9-1 downto 0);
signal st6col51: std_logic_vector(9-1 downto 0);
signal st6col52: std_logic_vector(8-1 downto 0);
signal st6col53: std_logic_vector(8-1 downto 0);
signal st6col54: std_logic_vector(7-1 downto 0);
signal st6col55: std_logic_vector(7-1 downto 0);
signal st6col56: std_logic_vector(6-1 downto 0);
signal st6col57: std_logic_vector(6-1 downto 0);
signal st6col58: std_logic_vector(5-1 downto 0);
signal st6col59: std_logic_vector(5-1 downto 0);
signal st6col60: std_logic_vector(4-1 downto 0);
signal st6col61: std_logic_vector(4-1 downto 0);
signal st6col62: std_logic_vector(3-1 downto 0);
signal st6col63: std_logic_vector(3-1 downto 0);
signal st6col64: std_logic_vector(2-1 downto 0);
signal st7col1: std_logic_vector(2-1 downto 0);
signal st7col2: std_logic_vector(1-1 downto 0);
signal st7col3: std_logic_vector(3-1 downto 0);
signal st7col4: std_logic_vector(2-1 downto 0);
signal st7col5: std_logic_vector(4-1 downto 0);
signal st7col6: std_logic_vector(3-1 downto 0);
signal st7col7: std_logic_vector(5-1 downto 0);
signal st7col8: std_logic_vector(4-1 downto 0);
signal st7col9: std_logic_vector(6-1 downto 0);
signal st7col10: std_logic_vector(5-1 downto 0);
signal st7col11: std_logic_vector(7-1 downto 0);
signal st7col12: std_logic_vector(6-1 downto 0);
signal st7col13: std_logic_vector(8-1 downto 0);
signal st7col14: std_logic_vector(7-1 downto 0);
signal st7col15: std_logic_vector(9-1 downto 0);
signal st7col16: std_logic_vector(8-1 downto 0);
signal st7col17: std_logic_vector(10-1 downto 0);
signal st7col18: std_logic_vector(9-1 downto 0);
signal st7col19: std_logic_vector(11-1 downto 0);
signal st7col20: std_logic_vector(10-1 downto 0);
signal st7col21: std_logic_vector(12-1 downto 0);
signal st7col22: std_logic_vector(11-1 downto 0);
signal st7col23: std_logic_vector(13-1 downto 0);
signal st7col24: std_logic_vector(12-1 downto 0);
signal st7col25: std_logic_vector(14-1 downto 0);
signal st7col26: std_logic_vector(13-1 downto 0);
signal st7col27: std_logic_vector(15-1 downto 0);
signal st7col28: std_logic_vector(14-1 downto 0);
signal st7col29: std_logic_vector(16-1 downto 0);
signal st7col30: std_logic_vector(15-1 downto 0);
signal st7col31: std_logic_vector(17-1 downto 0);
signal st7col32: std_logic_vector(16-1 downto 0);
signal st7col33: std_logic_vector(17-1 downto 0);
signal st7col34: std_logic_vector(17-1 downto 0);
signal st7col35: std_logic_vector(17-1 downto 0);
signal st7col36: std_logic_vector(17-1 downto 0);
signal st7col37: std_logic_vector(16-1 downto 0);
signal st7col38: std_logic_vector(15-1 downto 0);
signal st7col39: std_logic_vector(15-1 downto 0);
signal st7col40: std_logic_vector(14-1 downto 0);
signal st7col41: std_logic_vector(14-1 downto 0);
signal st7col42: std_logic_vector(13-1 downto 0);
signal st7col43: std_logic_vector(13-1 downto 0);
signal st7col44: std_logic_vector(12-1 downto 0);
signal st7col45: std_logic_vector(12-1 downto 0);
signal st7col46: std_logic_vector(11-1 downto 0);
signal st7col47: std_logic_vector(11-1 downto 0);
signal st7col48: std_logic_vector(10-1 downto 0);
signal st7col49: std_logic_vector(10-1 downto 0);
signal st7col50: std_logic_vector(9-1 downto 0);
signal st7col51: std_logic_vector(9-1 downto 0);
signal st7col52: std_logic_vector(8-1 downto 0);
signal st7col53: std_logic_vector(8-1 downto 0);
signal st7col54: std_logic_vector(7-1 downto 0);
signal st7col55: std_logic_vector(7-1 downto 0);
signal st7col56: std_logic_vector(6-1 downto 0);
signal st7col57: std_logic_vector(6-1 downto 0);
signal st7col58: std_logic_vector(5-1 downto 0);
signal st7col59: std_logic_vector(5-1 downto 0);
signal st7col60: std_logic_vector(4-1 downto 0);
signal st7col61: std_logic_vector(4-1 downto 0);
signal st7col62: std_logic_vector(3-1 downto 0);
signal st7col63: std_logic_vector(3-1 downto 0);
signal st7col64: std_logic_vector(2-1 downto 0);

-- END AUTOGEN DECL

begin
-- Extend multiplicand
a <= '0' & m_and;
a_neg_proc: process (a)
			begin
				for i in a'range loop
					a_neg(i) <= not a(i);
				end loop;
			end process;
			
a2_neg_proc: process (a2)
			begin
				for i in a2'range loop
					a2_neg(i) <= not a2(i);
				end loop;
			end process;
			
-- a2 = multiplicand * 2
a2 <= m_and & '0';

benc_proc: process(a, a2, a_neg, a2_neg, m_and, m_ier)
variable window: std_logic_vector(2 downto 0);
begin
	for i in 0 to N/2 loop
		if i = 0 then
			window := m_ier(1 downto 0) & '0';
		elsif i = N/2 then
			window := "00" & m_ier(N-1);
		else
			window := m_ier(2*i+1 downto 2*i-1);
		end if;
		
		if window = "000" then
			pprod(i) <= (OTHERS => '0');
		elsif window = "001" or window = "010" then
			pprod(i) <= a;
		elsif window = "101" or window = "110" then
			pprod(i) <= a_neg;
		elsif window = "011" then
			pprod(i) <= a2;
		elsif window = "100" then
			pprod(i) <= a2_neg;
		elsif window = "111" then
			pprod(i) <= (OTHERS => '1');
		end if;
		
	S(i) <= window(2);
	end loop;
end process;

-- BEGIN AUTOGEN COMPS
st6col1(0)<=st7col1(0);
st6col1(1)<=st7col1(1);
st6col2(0)<=st7col2(0);
st6col3(0)<=st7col3(0);
st6col3(1)<=st7col3(1);
st6col3(2)<=st7col3(2);
st6col4(0)<=st7col4(0);
st6col4(1)<=st7col4(1);
st6col5(0)<=st7col5(0);
st6col5(1)<=st7col5(1);
st6col5(2)<=st7col5(2);
st6col5(3)<=st7col5(3);
st6col6(0)<=st7col6(0);
st6col6(1)<=st7col6(1);
st6col6(2)<=st7col6(2);
st6col7(0)<=st7col7(0);
st6col7(1)<=st7col7(1);
st6col7(2)<=st7col7(2);
st6col7(3)<=st7col7(3);
st6col7(4)<=st7col7(4);
st6col8(0)<=st7col8(0);
st6col8(1)<=st7col8(1);
st6col8(2)<=st7col8(2);
st6col8(3)<=st7col8(3);
st6col9(0)<=st7col9(0);
st6col9(1)<=st7col9(1);
st6col9(2)<=st7col9(2);
st6col9(3)<=st7col9(3);
st6col9(4)<=st7col9(4);
st6col9(5)<=st7col9(5);
st6col10(0)<=st7col10(0);
st6col10(1)<=st7col10(1);
st6col10(2)<=st7col10(2);
st6col10(3)<=st7col10(3);
st6col10(4)<=st7col10(4);
st6col11(0)<=st7col11(0);
st6col11(1)<=st7col11(1);
st6col11(2)<=st7col11(2);
st6col11(3)<=st7col11(3);
st6col11(4)<=st7col11(4);
st6col11(5)<=st7col11(5);
st6col11(6)<=st7col11(6);
st6col12(0)<=st7col12(0);
st6col12(1)<=st7col12(1);
st6col12(2)<=st7col12(2);
st6col12(3)<=st7col12(3);
st6col12(4)<=st7col12(4);
st6col12(5)<=st7col12(5);
st6col13(0)<=st7col13(0);
st6col13(1)<=st7col13(1);
st6col13(2)<=st7col13(2);
st6col13(3)<=st7col13(3);
st6col13(4)<=st7col13(4);
st6col13(5)<=st7col13(5);
st6col13(6)<=st7col13(6);
st6col13(7)<=st7col13(7);
st6col14(0)<=st7col14(0);
st6col14(1)<=st7col14(1);
st6col14(2)<=st7col14(2);
st6col14(3)<=st7col14(3);
st6col14(4)<=st7col14(4);
st6col14(5)<=st7col14(5);
st6col14(6)<=st7col14(6);
st6col15(0)<=st7col15(0);
st6col15(1)<=st7col15(1);
st6col15(2)<=st7col15(2);
st6col15(3)<=st7col15(3);
st6col15(4)<=st7col15(4);
st6col15(5)<=st7col15(5);
st6col15(6)<=st7col15(6);
st6col15(7)<=st7col15(7);
st6col15(8)<=st7col15(8);
st6col16(0)<=st7col16(0);
st6col16(1)<=st7col16(1);
st6col16(2)<=st7col16(2);
st6col16(3)<=st7col16(3);
st6col16(4)<=st7col16(4);
st6col16(5)<=st7col16(5);
st6col16(6)<=st7col16(6);
st6col16(7)<=st7col16(7);
st6col17(0)<=st7col17(0);
st6col17(1)<=st7col17(1);
st6col17(2)<=st7col17(2);
st6col17(3)<=st7col17(3);
st6col17(4)<=st7col17(4);
st6col17(5)<=st7col17(5);
st6col17(6)<=st7col17(6);
st6col17(7)<=st7col17(7);
st6col17(8)<=st7col17(8);
st6col17(9)<=st7col17(9);
st6col18(0)<=st7col18(0);
st6col18(1)<=st7col18(1);
st6col18(2)<=st7col18(2);
st6col18(3)<=st7col18(3);
st6col18(4)<=st7col18(4);
st6col18(5)<=st7col18(5);
st6col18(6)<=st7col18(6);
st6col18(7)<=st7col18(7);
st6col18(8)<=st7col18(8);
st6col19(0)<=st7col19(0);
st6col19(1)<=st7col19(1);
st6col19(2)<=st7col19(2);
st6col19(3)<=st7col19(3);
st6col19(4)<=st7col19(4);
st6col19(5)<=st7col19(5);
st6col19(6)<=st7col19(6);
st6col19(7)<=st7col19(7);
st6col19(8)<=st7col19(8);
st6col19(9)<=st7col19(9);
st6col19(10)<=st7col19(10);
st6col20(0)<=st7col20(0);
st6col20(1)<=st7col20(1);
st6col20(2)<=st7col20(2);
st6col20(3)<=st7col20(3);
st6col20(4)<=st7col20(4);
st6col20(5)<=st7col20(5);
st6col20(6)<=st7col20(6);
st6col20(7)<=st7col20(7);
st6col20(8)<=st7col20(8);
st6col20(9)<=st7col20(9);
st6col21(0)<=st7col21(0);
st6col21(1)<=st7col21(1);
st6col21(2)<=st7col21(2);
st6col21(3)<=st7col21(3);
st6col21(4)<=st7col21(4);
st6col21(5)<=st7col21(5);
st6col21(6)<=st7col21(6);
st6col21(7)<=st7col21(7);
st6col21(8)<=st7col21(8);
st6col21(9)<=st7col21(9);
st6col21(10)<=st7col21(10);
st6col21(11)<=st7col21(11);
st6col22(0)<=st7col22(0);
st6col22(1)<=st7col22(1);
st6col22(2)<=st7col22(2);
st6col22(3)<=st7col22(3);
st6col22(4)<=st7col22(4);
st6col22(5)<=st7col22(5);
st6col22(6)<=st7col22(6);
st6col22(7)<=st7col22(7);
st6col22(8)<=st7col22(8);
st6col22(9)<=st7col22(9);
st6col22(10)<=st7col22(10);
st6col23(0)<=st7col23(0);
st6col23(1)<=st7col23(1);
st6col23(2)<=st7col23(2);
st6col23(3)<=st7col23(3);
st6col23(4)<=st7col23(4);
st6col23(5)<=st7col23(5);
st6col23(6)<=st7col23(6);
st6col23(7)<=st7col23(7);
st6col23(8)<=st7col23(8);
st6col23(9)<=st7col23(9);
st6col23(10)<=st7col23(10);
st6col23(11)<=st7col23(11);
st6col23(12)<=st7col23(12);
st6col24(0)<=st7col24(0);
st6col24(1)<=st7col24(1);
st6col24(2)<=st7col24(2);
st6col24(3)<=st7col24(3);
st6col24(4)<=st7col24(4);
st6col24(5)<=st7col24(5);
st6col24(6)<=st7col24(6);
st6col24(7)<=st7col24(7);
st6col24(8)<=st7col24(8);
st6col24(9)<=st7col24(9);
st6col24(10)<=st7col24(10);
st6col24(11)<=st7col24(11);
ha1st7col25: HA port map(st7col25(0),st7col25(1),st6col25(0),st6col26(0));
st6col25(1)<=st7col25(2);
st6col25(2)<=st7col25(3);
st6col25(3)<=st7col25(4);
st6col25(4)<=st7col25(5);
st6col25(5)<=st7col25(6);
st6col25(6)<=st7col25(7);
st6col25(7)<=st7col25(8);
st6col25(8)<=st7col25(9);
st6col25(9)<=st7col25(10);
st6col25(10)<=st7col25(11);
st6col25(11)<=st7col25(12);
st6col25(12)<=st7col25(13);
ha1st7col26: HA port map(st7col26(0),st7col26(1),st6col26(1),st6col27(0));
st6col26(2)<=st7col26(2);
st6col26(3)<=st7col26(3);
st6col26(4)<=st7col26(4);
st6col26(5)<=st7col26(5);
st6col26(6)<=st7col26(6);
st6col26(7)<=st7col26(7);
st6col26(8)<=st7col26(8);
st6col26(9)<=st7col26(9);
st6col26(10)<=st7col26(10);
st6col26(11)<=st7col26(11);
st6col26(12)<=st7col26(12);
fa0st7col27: FA port map(st7col27(0),st7col27(1),st7col27(2),st6col27(1),st6col28(0));
ha1st7col27: HA port map(st7col27(3),st7col27(4),st6col27(2),st6col28(1));
st6col27(3)<=st7col27(5);
st6col27(4)<=st7col27(6);
st6col27(5)<=st7col27(7);
st6col27(6)<=st7col27(8);
st6col27(7)<=st7col27(9);
st6col27(8)<=st7col27(10);
st6col27(9)<=st7col27(11);
st6col27(10)<=st7col27(12);
st6col27(11)<=st7col27(13);
st6col27(12)<=st7col27(14);
fa0st7col28: FA port map(st7col28(0),st7col28(1),st7col28(2),st6col28(2),st6col29(0));
ha1st7col28: HA port map(st7col28(3),st7col28(4),st6col28(3),st6col29(1));
st6col28(4)<=st7col28(5);
st6col28(5)<=st7col28(6);
st6col28(6)<=st7col28(7);
st6col28(7)<=st7col28(8);
st6col28(8)<=st7col28(9);
st6col28(9)<=st7col28(10);
st6col28(10)<=st7col28(11);
st6col28(11)<=st7col28(12);
st6col28(12)<=st7col28(13);
fa0st7col29: FA port map(st7col29(0),st7col29(1),st7col29(2),st6col29(2),st6col30(0));
fa1st7col29: FA port map(st7col29(3),st7col29(4),st7col29(5),st6col29(3),st6col30(1));
ha1st7col29: HA port map(st7col29(6),st7col29(7),st6col29(4),st6col30(2));
st6col29(5)<=st7col29(8);
st6col29(6)<=st7col29(9);
st6col29(7)<=st7col29(10);
st6col29(8)<=st7col29(11);
st6col29(9)<=st7col29(12);
st6col29(10)<=st7col29(13);
st6col29(11)<=st7col29(14);
st6col29(12)<=st7col29(15);
fa0st7col30: FA port map(st7col30(0),st7col30(1),st7col30(2),st6col30(3),st6col31(0));
fa1st7col30: FA port map(st7col30(3),st7col30(4),st7col30(5),st6col30(4),st6col31(1));
ha1st7col30: HA port map(st7col30(6),st7col30(7),st6col30(5),st6col31(2));
st6col30(6)<=st7col30(8);
st6col30(7)<=st7col30(9);
st6col30(8)<=st7col30(10);
st6col30(9)<=st7col30(11);
st6col30(10)<=st7col30(12);
st6col30(11)<=st7col30(13);
st6col30(12)<=st7col30(14);
fa0st7col31: FA port map(st7col31(0),st7col31(1),st7col31(2),st6col31(3),st6col32(0));
fa1st7col31: FA port map(st7col31(3),st7col31(4),st7col31(5),st6col31(4),st6col32(1));
fa2st7col31: FA port map(st7col31(6),st7col31(7),st7col31(8),st6col31(5),st6col32(2));
ha1st7col31: HA port map(st7col31(9),st7col31(10),st6col31(6),st6col32(3));
st6col31(7)<=st7col31(11);
st6col31(8)<=st7col31(12);
st6col31(9)<=st7col31(13);
st6col31(10)<=st7col31(14);
st6col31(11)<=st7col31(15);
st6col31(12)<=st7col31(16);
fa0st7col32: FA port map(st7col32(0),st7col32(1),st7col32(2),st6col32(4),st6col33(0));
fa1st7col32: FA port map(st7col32(3),st7col32(4),st7col32(5),st6col32(5),st6col33(1));
fa2st7col32: FA port map(st7col32(6),st7col32(7),st7col32(8),st6col32(6),st6col33(2));
ha1st7col32: HA port map(st7col32(9),st7col32(10),st6col32(7),st6col33(3));
st6col32(8)<=st7col32(11);
st6col32(9)<=st7col32(12);
st6col32(10)<=st7col32(13);
st6col32(11)<=st7col32(14);
st6col32(12)<=st7col32(15);
fa0st7col33: FA port map(st7col33(0),st7col33(1),st7col33(2),st6col33(4),st6col34(0));
fa1st7col33: FA port map(st7col33(3),st7col33(4),st7col33(5),st6col33(5),st6col34(1));
fa2st7col33: FA port map(st7col33(6),st7col33(7),st7col33(8),st6col33(6),st6col34(2));
fa3st7col33: FA port map(st7col33(9),st7col33(10),st7col33(11),st6col33(7),st6col34(3));
st6col33(8)<=st7col33(12);
st6col33(9)<=st7col33(13);
st6col33(10)<=st7col33(14);
st6col33(11)<=st7col33(15);
st6col33(12)<=st7col33(16);
fa0st7col34: FA port map(st7col34(0),st7col34(1),st7col34(2),st6col34(4),st6col35(0));
fa1st7col34: FA port map(st7col34(3),st7col34(4),st7col34(5),st6col34(5),st6col35(1));
fa2st7col34: FA port map(st7col34(6),st7col34(7),st7col34(8),st6col34(6),st6col35(2));
fa3st7col34: FA port map(st7col34(9),st7col34(10),st7col34(11),st6col34(7),st6col35(3));
st6col34(8)<=st7col34(12);
st6col34(9)<=st7col34(13);
st6col34(10)<=st7col34(14);
st6col34(11)<=st7col34(15);
st6col34(12)<=st7col34(16);
fa0st7col35: FA port map(st7col35(0),st7col35(1),st7col35(2),st6col35(4),st6col36(0));
fa1st7col35: FA port map(st7col35(3),st7col35(4),st7col35(5),st6col35(5),st6col36(1));
fa2st7col35: FA port map(st7col35(6),st7col35(7),st7col35(8),st6col35(6),st6col36(2));
fa3st7col35: FA port map(st7col35(9),st7col35(10),st7col35(11),st6col35(7),st6col36(3));
st6col35(8)<=st7col35(12);
st6col35(9)<=st7col35(13);
st6col35(10)<=st7col35(14);
st6col35(11)<=st7col35(15);
st6col35(12)<=st7col35(16);
fa0st7col36: FA port map(st7col36(0),st7col36(1),st7col36(2),st6col36(4),st6col37(0));
fa1st7col36: FA port map(st7col36(3),st7col36(4),st7col36(5),st6col36(5),st6col37(1));
fa2st7col36: FA port map(st7col36(6),st7col36(7),st7col36(8),st6col36(6),st6col37(2));
fa3st7col36: FA port map(st7col36(9),st7col36(10),st7col36(11),st6col36(7),st6col37(3));
st6col36(8)<=st7col36(12);
st6col36(9)<=st7col36(13);
st6col36(10)<=st7col36(14);
st6col36(11)<=st7col36(15);
st6col36(12)<=st7col36(16);
fa0st7col37: FA port map(st7col37(0),st7col37(1),st7col37(2),st6col37(4),st6col38(0));
fa1st7col37: FA port map(st7col37(3),st7col37(4),st7col37(5),st6col37(5),st6col38(1));
fa2st7col37: FA port map(st7col37(6),st7col37(7),st7col37(8),st6col37(6),st6col38(2));
ha1st7col37: HA port map(st7col37(9),st7col37(10),st6col37(7),st6col38(3));
st6col37(8)<=st7col37(11);
st6col37(9)<=st7col37(12);
st6col37(10)<=st7col37(13);
st6col37(11)<=st7col37(14);
st6col37(12)<=st7col37(15);
fa0st7col38: FA port map(st7col38(0),st7col38(1),st7col38(2),st6col38(4),st6col39(0));
fa1st7col38: FA port map(st7col38(3),st7col38(4),st7col38(5),st6col38(5),st6col39(1));
fa2st7col38: FA port map(st7col38(6),st7col38(7),st7col38(8),st6col38(6),st6col39(2));
st6col38(7)<=st7col38(9);
st6col38(8)<=st7col38(10);
st6col38(9)<=st7col38(11);
st6col38(10)<=st7col38(12);
st6col38(11)<=st7col38(13);
st6col38(12)<=st7col38(14);
fa0st7col39: FA port map(st7col39(0),st7col39(1),st7col39(2),st6col39(3),st6col40(0));
fa1st7col39: FA port map(st7col39(3),st7col39(4),st7col39(5),st6col39(4),st6col40(1));
ha1st7col39: HA port map(st7col39(6),st7col39(7),st6col39(5),st6col40(2));
st6col39(6)<=st7col39(8);
st6col39(7)<=st7col39(9);
st6col39(8)<=st7col39(10);
st6col39(9)<=st7col39(11);
st6col39(10)<=st7col39(12);
st6col39(11)<=st7col39(13);
st6col39(12)<=st7col39(14);
fa0st7col40: FA port map(st7col40(0),st7col40(1),st7col40(2),st6col40(3),st6col41(0));
fa1st7col40: FA port map(st7col40(3),st7col40(4),st7col40(5),st6col40(4),st6col41(1));
st6col40(5)<=st7col40(6);
st6col40(6)<=st7col40(7);
st6col40(7)<=st7col40(8);
st6col40(8)<=st7col40(9);
st6col40(9)<=st7col40(10);
st6col40(10)<=st7col40(11);
st6col40(11)<=st7col40(12);
st6col40(12)<=st7col40(13);
fa0st7col41: FA port map(st7col41(0),st7col41(1),st7col41(2),st6col41(2),st6col42(0));
ha1st7col41: HA port map(st7col41(3),st7col41(4),st6col41(3),st6col42(1));
st6col41(4)<=st7col41(5);
st6col41(5)<=st7col41(6);
st6col41(6)<=st7col41(7);
st6col41(7)<=st7col41(8);
st6col41(8)<=st7col41(9);
st6col41(9)<=st7col41(10);
st6col41(10)<=st7col41(11);
st6col41(11)<=st7col41(12);
st6col41(12)<=st7col41(13);
fa0st7col42: FA port map(st7col42(0),st7col42(1),st7col42(2),st6col42(2),st6col43(0));
st6col42(3)<=st7col42(3);
st6col42(4)<=st7col42(4);
st6col42(5)<=st7col42(5);
st6col42(6)<=st7col42(6);
st6col42(7)<=st7col42(7);
st6col42(8)<=st7col42(8);
st6col42(9)<=st7col42(9);
st6col42(10)<=st7col42(10);
st6col42(11)<=st7col42(11);
st6col42(12)<=st7col42(12);
ha1st7col43: HA port map(st7col43(0),st7col43(1),st6col43(1),st6col44(0));
st6col43(2)<=st7col43(2);
st6col43(3)<=st7col43(3);
st6col43(4)<=st7col43(4);
st6col43(5)<=st7col43(5);
st6col43(6)<=st7col43(6);
st6col43(7)<=st7col43(7);
st6col43(8)<=st7col43(8);
st6col43(9)<=st7col43(9);
st6col43(10)<=st7col43(10);
st6col43(11)<=st7col43(11);
st6col43(12)<=st7col43(12);
st6col44(1)<=st7col44(0);
st6col44(2)<=st7col44(1);
st6col44(3)<=st7col44(2);
st6col44(4)<=st7col44(3);
st6col44(5)<=st7col44(4);
st6col44(6)<=st7col44(5);
st6col44(7)<=st7col44(6);
st6col44(8)<=st7col44(7);
st6col44(9)<=st7col44(8);
st6col44(10)<=st7col44(9);
st6col44(11)<=st7col44(10);
st6col44(12)<=st7col44(11);
st6col45(0)<=st7col45(0);
st6col45(1)<=st7col45(1);
st6col45(2)<=st7col45(2);
st6col45(3)<=st7col45(3);
st6col45(4)<=st7col45(4);
st6col45(5)<=st7col45(5);
st6col45(6)<=st7col45(6);
st6col45(7)<=st7col45(7);
st6col45(8)<=st7col45(8);
st6col45(9)<=st7col45(9);
st6col45(10)<=st7col45(10);
st6col45(11)<=st7col45(11);
st6col46(0)<=st7col46(0);
st6col46(1)<=st7col46(1);
st6col46(2)<=st7col46(2);
st6col46(3)<=st7col46(3);
st6col46(4)<=st7col46(4);
st6col46(5)<=st7col46(5);
st6col46(6)<=st7col46(6);
st6col46(7)<=st7col46(7);
st6col46(8)<=st7col46(8);
st6col46(9)<=st7col46(9);
st6col46(10)<=st7col46(10);
st6col47(0)<=st7col47(0);
st6col47(1)<=st7col47(1);
st6col47(2)<=st7col47(2);
st6col47(3)<=st7col47(3);
st6col47(4)<=st7col47(4);
st6col47(5)<=st7col47(5);
st6col47(6)<=st7col47(6);
st6col47(7)<=st7col47(7);
st6col47(8)<=st7col47(8);
st6col47(9)<=st7col47(9);
st6col47(10)<=st7col47(10);
st6col48(0)<=st7col48(0);
st6col48(1)<=st7col48(1);
st6col48(2)<=st7col48(2);
st6col48(3)<=st7col48(3);
st6col48(4)<=st7col48(4);
st6col48(5)<=st7col48(5);
st6col48(6)<=st7col48(6);
st6col48(7)<=st7col48(7);
st6col48(8)<=st7col48(8);
st6col48(9)<=st7col48(9);
st6col49(0)<=st7col49(0);
st6col49(1)<=st7col49(1);
st6col49(2)<=st7col49(2);
st6col49(3)<=st7col49(3);
st6col49(4)<=st7col49(4);
st6col49(5)<=st7col49(5);
st6col49(6)<=st7col49(6);
st6col49(7)<=st7col49(7);
st6col49(8)<=st7col49(8);
st6col49(9)<=st7col49(9);
st6col50(0)<=st7col50(0);
st6col50(1)<=st7col50(1);
st6col50(2)<=st7col50(2);
st6col50(3)<=st7col50(3);
st6col50(4)<=st7col50(4);
st6col50(5)<=st7col50(5);
st6col50(6)<=st7col50(6);
st6col50(7)<=st7col50(7);
st6col50(8)<=st7col50(8);
st6col51(0)<=st7col51(0);
st6col51(1)<=st7col51(1);
st6col51(2)<=st7col51(2);
st6col51(3)<=st7col51(3);
st6col51(4)<=st7col51(4);
st6col51(5)<=st7col51(5);
st6col51(6)<=st7col51(6);
st6col51(7)<=st7col51(7);
st6col51(8)<=st7col51(8);
st6col52(0)<=st7col52(0);
st6col52(1)<=st7col52(1);
st6col52(2)<=st7col52(2);
st6col52(3)<=st7col52(3);
st6col52(4)<=st7col52(4);
st6col52(5)<=st7col52(5);
st6col52(6)<=st7col52(6);
st6col52(7)<=st7col52(7);
st6col53(0)<=st7col53(0);
st6col53(1)<=st7col53(1);
st6col53(2)<=st7col53(2);
st6col53(3)<=st7col53(3);
st6col53(4)<=st7col53(4);
st6col53(5)<=st7col53(5);
st6col53(6)<=st7col53(6);
st6col53(7)<=st7col53(7);
st6col54(0)<=st7col54(0);
st6col54(1)<=st7col54(1);
st6col54(2)<=st7col54(2);
st6col54(3)<=st7col54(3);
st6col54(4)<=st7col54(4);
st6col54(5)<=st7col54(5);
st6col54(6)<=st7col54(6);
st6col55(0)<=st7col55(0);
st6col55(1)<=st7col55(1);
st6col55(2)<=st7col55(2);
st6col55(3)<=st7col55(3);
st6col55(4)<=st7col55(4);
st6col55(5)<=st7col55(5);
st6col55(6)<=st7col55(6);
st6col56(0)<=st7col56(0);
st6col56(1)<=st7col56(1);
st6col56(2)<=st7col56(2);
st6col56(3)<=st7col56(3);
st6col56(4)<=st7col56(4);
st6col56(5)<=st7col56(5);
st6col57(0)<=st7col57(0);
st6col57(1)<=st7col57(1);
st6col57(2)<=st7col57(2);
st6col57(3)<=st7col57(3);
st6col57(4)<=st7col57(4);
st6col57(5)<=st7col57(5);
st6col58(0)<=st7col58(0);
st6col58(1)<=st7col58(1);
st6col58(2)<=st7col58(2);
st6col58(3)<=st7col58(3);
st6col58(4)<=st7col58(4);
st6col59(0)<=st7col59(0);
st6col59(1)<=st7col59(1);
st6col59(2)<=st7col59(2);
st6col59(3)<=st7col59(3);
st6col59(4)<=st7col59(4);
st6col60(0)<=st7col60(0);
st6col60(1)<=st7col60(1);
st6col60(2)<=st7col60(2);
st6col60(3)<=st7col60(3);
st6col61(0)<=st7col61(0);
st6col61(1)<=st7col61(1);
st6col61(2)<=st7col61(2);
st6col61(3)<=st7col61(3);
st6col62(0)<=st7col62(0);
st6col62(1)<=st7col62(1);
st6col62(2)<=st7col62(2);
st6col63(0)<=st7col63(0);
st6col63(1)<=st7col63(1);
st6col63(2)<=st7col63(2);
st6col64(0)<=st7col64(0);
st6col64(1)<=st7col64(1);
st5col1(0)<=st6col1(0);
st5col1(1)<=st6col1(1);
st5col2(0)<=st6col2(0);
st5col3(0)<=st6col3(0);
st5col3(1)<=st6col3(1);
st5col3(2)<=st6col3(2);
st5col4(0)<=st6col4(0);
st5col4(1)<=st6col4(1);
st5col5(0)<=st6col5(0);
st5col5(1)<=st6col5(1);
st5col5(2)<=st6col5(2);
st5col5(3)<=st6col5(3);
st5col6(0)<=st6col6(0);
st5col6(1)<=st6col6(1);
st5col6(2)<=st6col6(2);
st5col7(0)<=st6col7(0);
st5col7(1)<=st6col7(1);
st5col7(2)<=st6col7(2);
st5col7(3)<=st6col7(3);
st5col7(4)<=st6col7(4);
st5col8(0)<=st6col8(0);
st5col8(1)<=st6col8(1);
st5col8(2)<=st6col8(2);
st5col8(3)<=st6col8(3);
st5col9(0)<=st6col9(0);
st5col9(1)<=st6col9(1);
st5col9(2)<=st6col9(2);
st5col9(3)<=st6col9(3);
st5col9(4)<=st6col9(4);
st5col9(5)<=st6col9(5);
st5col10(0)<=st6col10(0);
st5col10(1)<=st6col10(1);
st5col10(2)<=st6col10(2);
st5col10(3)<=st6col10(3);
st5col10(4)<=st6col10(4);
st5col11(0)<=st6col11(0);
st5col11(1)<=st6col11(1);
st5col11(2)<=st6col11(2);
st5col11(3)<=st6col11(3);
st5col11(4)<=st6col11(4);
st5col11(5)<=st6col11(5);
st5col11(6)<=st6col11(6);
st5col12(0)<=st6col12(0);
st5col12(1)<=st6col12(1);
st5col12(2)<=st6col12(2);
st5col12(3)<=st6col12(3);
st5col12(4)<=st6col12(4);
st5col12(5)<=st6col12(5);
st5col13(0)<=st6col13(0);
st5col13(1)<=st6col13(1);
st5col13(2)<=st6col13(2);
st5col13(3)<=st6col13(3);
st5col13(4)<=st6col13(4);
st5col13(5)<=st6col13(5);
st5col13(6)<=st6col13(6);
st5col13(7)<=st6col13(7);
st5col14(0)<=st6col14(0);
st5col14(1)<=st6col14(1);
st5col14(2)<=st6col14(2);
st5col14(3)<=st6col14(3);
st5col14(4)<=st6col14(4);
st5col14(5)<=st6col14(5);
st5col14(6)<=st6col14(6);
st5col15(0)<=st6col15(0);
st5col15(1)<=st6col15(1);
st5col15(2)<=st6col15(2);
st5col15(3)<=st6col15(3);
st5col15(4)<=st6col15(4);
st5col15(5)<=st6col15(5);
st5col15(6)<=st6col15(6);
st5col15(7)<=st6col15(7);
st5col15(8)<=st6col15(8);
st5col16(0)<=st6col16(0);
st5col16(1)<=st6col16(1);
st5col16(2)<=st6col16(2);
st5col16(3)<=st6col16(3);
st5col16(4)<=st6col16(4);
st5col16(5)<=st6col16(5);
st5col16(6)<=st6col16(6);
st5col16(7)<=st6col16(7);
ha1st6col17: HA port map(st6col17(0),st6col17(1),st5col17(0),st5col18(0));
st5col17(1)<=st6col17(2);
st5col17(2)<=st6col17(3);
st5col17(3)<=st6col17(4);
st5col17(4)<=st6col17(5);
st5col17(5)<=st6col17(6);
st5col17(6)<=st6col17(7);
st5col17(7)<=st6col17(8);
st5col17(8)<=st6col17(9);
ha1st6col18: HA port map(st6col18(0),st6col18(1),st5col18(1),st5col19(0));
st5col18(2)<=st6col18(2);
st5col18(3)<=st6col18(3);
st5col18(4)<=st6col18(4);
st5col18(5)<=st6col18(5);
st5col18(6)<=st6col18(6);
st5col18(7)<=st6col18(7);
st5col18(8)<=st6col18(8);
fa0st6col19: FA port map(st6col19(0),st6col19(1),st6col19(2),st5col19(1),st5col20(0));
ha1st6col19: HA port map(st6col19(3),st6col19(4),st5col19(2),st5col20(1));
st5col19(3)<=st6col19(5);
st5col19(4)<=st6col19(6);
st5col19(5)<=st6col19(7);
st5col19(6)<=st6col19(8);
st5col19(7)<=st6col19(9);
st5col19(8)<=st6col19(10);
fa0st6col20: FA port map(st6col20(0),st6col20(1),st6col20(2),st5col20(2),st5col21(0));
ha1st6col20: HA port map(st6col20(3),st6col20(4),st5col20(3),st5col21(1));
st5col20(4)<=st6col20(5);
st5col20(5)<=st6col20(6);
st5col20(6)<=st6col20(7);
st5col20(7)<=st6col20(8);
st5col20(8)<=st6col20(9);
fa0st6col21: FA port map(st6col21(0),st6col21(1),st6col21(2),st5col21(2),st5col22(0));
fa1st6col21: FA port map(st6col21(3),st6col21(4),st6col21(5),st5col21(3),st5col22(1));
ha1st6col21: HA port map(st6col21(6),st6col21(7),st5col21(4),st5col22(2));
st5col21(5)<=st6col21(8);
st5col21(6)<=st6col21(9);
st5col21(7)<=st6col21(10);
st5col21(8)<=st6col21(11);
fa0st6col22: FA port map(st6col22(0),st6col22(1),st6col22(2),st5col22(3),st5col23(0));
fa1st6col22: FA port map(st6col22(3),st6col22(4),st6col22(5),st5col22(4),st5col23(1));
ha1st6col22: HA port map(st6col22(6),st6col22(7),st5col22(5),st5col23(2));
st5col22(6)<=st6col22(8);
st5col22(7)<=st6col22(9);
st5col22(8)<=st6col22(10);
fa0st6col23: FA port map(st6col23(0),st6col23(1),st6col23(2),st5col23(3),st5col24(0));
fa1st6col23: FA port map(st6col23(3),st6col23(4),st6col23(5),st5col23(4),st5col24(1));
fa2st6col23: FA port map(st6col23(6),st6col23(7),st6col23(8),st5col23(5),st5col24(2));
ha1st6col23: HA port map(st6col23(9),st6col23(10),st5col23(6),st5col24(3));
st5col23(7)<=st6col23(11);
st5col23(8)<=st6col23(12);
fa0st6col24: FA port map(st6col24(0),st6col24(1),st6col24(2),st5col24(4),st5col25(0));
fa1st6col24: FA port map(st6col24(3),st6col24(4),st6col24(5),st5col24(5),st5col25(1));
fa2st6col24: FA port map(st6col24(6),st6col24(7),st6col24(8),st5col24(6),st5col25(2));
ha1st6col24: HA port map(st6col24(9),st6col24(10),st5col24(7),st5col25(3));
st5col24(8)<=st6col24(11);
fa0st6col25: FA port map(st6col25(0),st6col25(1),st6col25(2),st5col25(4),st5col26(0));
fa1st6col25: FA port map(st6col25(3),st6col25(4),st6col25(5),st5col25(5),st5col26(1));
fa2st6col25: FA port map(st6col25(6),st6col25(7),st6col25(8),st5col25(6),st5col26(2));
fa3st6col25: FA port map(st6col25(9),st6col25(10),st6col25(11),st5col25(7),st5col26(3));
st5col25(8)<=st6col25(12);
fa0st6col26: FA port map(st6col26(0),st6col26(1),st6col26(2),st5col26(4),st5col27(0));
fa1st6col26: FA port map(st6col26(3),st6col26(4),st6col26(5),st5col26(5),st5col27(1));
fa2st6col26: FA port map(st6col26(6),st6col26(7),st6col26(8),st5col26(6),st5col27(2));
fa3st6col26: FA port map(st6col26(9),st6col26(10),st6col26(11),st5col26(7),st5col27(3));
st5col26(8)<=st6col26(12);
fa0st6col27: FA port map(st6col27(0),st6col27(1),st6col27(2),st5col27(4),st5col28(0));
fa1st6col27: FA port map(st6col27(3),st6col27(4),st6col27(5),st5col27(5),st5col28(1));
fa2st6col27: FA port map(st6col27(6),st6col27(7),st6col27(8),st5col27(6),st5col28(2));
fa3st6col27: FA port map(st6col27(9),st6col27(10),st6col27(11),st5col27(7),st5col28(3));
st5col27(8)<=st6col27(12);
fa0st6col28: FA port map(st6col28(0),st6col28(1),st6col28(2),st5col28(4),st5col29(0));
fa1st6col28: FA port map(st6col28(3),st6col28(4),st6col28(5),st5col28(5),st5col29(1));
fa2st6col28: FA port map(st6col28(6),st6col28(7),st6col28(8),st5col28(6),st5col29(2));
fa3st6col28: FA port map(st6col28(9),st6col28(10),st6col28(11),st5col28(7),st5col29(3));
st5col28(8)<=st6col28(12);
fa0st6col29: FA port map(st6col29(0),st6col29(1),st6col29(2),st5col29(4),st5col30(0));
fa1st6col29: FA port map(st6col29(3),st6col29(4),st6col29(5),st5col29(5),st5col30(1));
fa2st6col29: FA port map(st6col29(6),st6col29(7),st6col29(8),st5col29(6),st5col30(2));
fa3st6col29: FA port map(st6col29(9),st6col29(10),st6col29(11),st5col29(7),st5col30(3));
st5col29(8)<=st6col29(12);
fa0st6col30: FA port map(st6col30(0),st6col30(1),st6col30(2),st5col30(4),st5col31(0));
fa1st6col30: FA port map(st6col30(3),st6col30(4),st6col30(5),st5col30(5),st5col31(1));
fa2st6col30: FA port map(st6col30(6),st6col30(7),st6col30(8),st5col30(6),st5col31(2));
fa3st6col30: FA port map(st6col30(9),st6col30(10),st6col30(11),st5col30(7),st5col31(3));
st5col30(8)<=st6col30(12);
fa0st6col31: FA port map(st6col31(0),st6col31(1),st6col31(2),st5col31(4),st5col32(0));
fa1st6col31: FA port map(st6col31(3),st6col31(4),st6col31(5),st5col31(5),st5col32(1));
fa2st6col31: FA port map(st6col31(6),st6col31(7),st6col31(8),st5col31(6),st5col32(2));
fa3st6col31: FA port map(st6col31(9),st6col31(10),st6col31(11),st5col31(7),st5col32(3));
st5col31(8)<=st6col31(12);
fa0st6col32: FA port map(st6col32(0),st6col32(1),st6col32(2),st5col32(4),st5col33(0));
fa1st6col32: FA port map(st6col32(3),st6col32(4),st6col32(5),st5col32(5),st5col33(1));
fa2st6col32: FA port map(st6col32(6),st6col32(7),st6col32(8),st5col32(6),st5col33(2));
fa3st6col32: FA port map(st6col32(9),st6col32(10),st6col32(11),st5col32(7),st5col33(3));
st5col32(8)<=st6col32(12);
fa0st6col33: FA port map(st6col33(0),st6col33(1),st6col33(2),st5col33(4),st5col34(0));
fa1st6col33: FA port map(st6col33(3),st6col33(4),st6col33(5),st5col33(5),st5col34(1));
fa2st6col33: FA port map(st6col33(6),st6col33(7),st6col33(8),st5col33(6),st5col34(2));
fa3st6col33: FA port map(st6col33(9),st6col33(10),st6col33(11),st5col33(7),st5col34(3));
st5col33(8)<=st6col33(12);
fa0st6col34: FA port map(st6col34(0),st6col34(1),st6col34(2),st5col34(4),st5col35(0));
fa1st6col34: FA port map(st6col34(3),st6col34(4),st6col34(5),st5col34(5),st5col35(1));
fa2st6col34: FA port map(st6col34(6),st6col34(7),st6col34(8),st5col34(6),st5col35(2));
fa3st6col34: FA port map(st6col34(9),st6col34(10),st6col34(11),st5col34(7),st5col35(3));
st5col34(8)<=st6col34(12);
fa0st6col35: FA port map(st6col35(0),st6col35(1),st6col35(2),st5col35(4),st5col36(0));
fa1st6col35: FA port map(st6col35(3),st6col35(4),st6col35(5),st5col35(5),st5col36(1));
fa2st6col35: FA port map(st6col35(6),st6col35(7),st6col35(8),st5col35(6),st5col36(2));
fa3st6col35: FA port map(st6col35(9),st6col35(10),st6col35(11),st5col35(7),st5col36(3));
st5col35(8)<=st6col35(12);
fa0st6col36: FA port map(st6col36(0),st6col36(1),st6col36(2),st5col36(4),st5col37(0));
fa1st6col36: FA port map(st6col36(3),st6col36(4),st6col36(5),st5col36(5),st5col37(1));
fa2st6col36: FA port map(st6col36(6),st6col36(7),st6col36(8),st5col36(6),st5col37(2));
fa3st6col36: FA port map(st6col36(9),st6col36(10),st6col36(11),st5col36(7),st5col37(3));
st5col36(8)<=st6col36(12);
fa0st6col37: FA port map(st6col37(0),st6col37(1),st6col37(2),st5col37(4),st5col38(0));
fa1st6col37: FA port map(st6col37(3),st6col37(4),st6col37(5),st5col37(5),st5col38(1));
fa2st6col37: FA port map(st6col37(6),st6col37(7),st6col37(8),st5col37(6),st5col38(2));
fa3st6col37: FA port map(st6col37(9),st6col37(10),st6col37(11),st5col37(7),st5col38(3));
st5col37(8)<=st6col37(12);
fa0st6col38: FA port map(st6col38(0),st6col38(1),st6col38(2),st5col38(4),st5col39(0));
fa1st6col38: FA port map(st6col38(3),st6col38(4),st6col38(5),st5col38(5),st5col39(1));
fa2st6col38: FA port map(st6col38(6),st6col38(7),st6col38(8),st5col38(6),st5col39(2));
fa3st6col38: FA port map(st6col38(9),st6col38(10),st6col38(11),st5col38(7),st5col39(3));
st5col38(8)<=st6col38(12);
fa0st6col39: FA port map(st6col39(0),st6col39(1),st6col39(2),st5col39(4),st5col40(0));
fa1st6col39: FA port map(st6col39(3),st6col39(4),st6col39(5),st5col39(5),st5col40(1));
fa2st6col39: FA port map(st6col39(6),st6col39(7),st6col39(8),st5col39(6),st5col40(2));
fa3st6col39: FA port map(st6col39(9),st6col39(10),st6col39(11),st5col39(7),st5col40(3));
st5col39(8)<=st6col39(12);
fa0st6col40: FA port map(st6col40(0),st6col40(1),st6col40(2),st5col40(4),st5col41(0));
fa1st6col40: FA port map(st6col40(3),st6col40(4),st6col40(5),st5col40(5),st5col41(1));
fa2st6col40: FA port map(st6col40(6),st6col40(7),st6col40(8),st5col40(6),st5col41(2));
fa3st6col40: FA port map(st6col40(9),st6col40(10),st6col40(11),st5col40(7),st5col41(3));
st5col40(8)<=st6col40(12);
fa0st6col41: FA port map(st6col41(0),st6col41(1),st6col41(2),st5col41(4),st5col42(0));
fa1st6col41: FA port map(st6col41(3),st6col41(4),st6col41(5),st5col41(5),st5col42(1));
fa2st6col41: FA port map(st6col41(6),st6col41(7),st6col41(8),st5col41(6),st5col42(2));
fa3st6col41: FA port map(st6col41(9),st6col41(10),st6col41(11),st5col41(7),st5col42(3));
st5col41(8)<=st6col41(12);
fa0st6col42: FA port map(st6col42(0),st6col42(1),st6col42(2),st5col42(4),st5col43(0));
fa1st6col42: FA port map(st6col42(3),st6col42(4),st6col42(5),st5col42(5),st5col43(1));
fa2st6col42: FA port map(st6col42(6),st6col42(7),st6col42(8),st5col42(6),st5col43(2));
fa3st6col42: FA port map(st6col42(9),st6col42(10),st6col42(11),st5col42(7),st5col43(3));
st5col42(8)<=st6col42(12);
fa0st6col43: FA port map(st6col43(0),st6col43(1),st6col43(2),st5col43(4),st5col44(0));
fa1st6col43: FA port map(st6col43(3),st6col43(4),st6col43(5),st5col43(5),st5col44(1));
fa2st6col43: FA port map(st6col43(6),st6col43(7),st6col43(8),st5col43(6),st5col44(2));
fa3st6col43: FA port map(st6col43(9),st6col43(10),st6col43(11),st5col43(7),st5col44(3));
st5col43(8)<=st6col43(12);
fa0st6col44: FA port map(st6col44(0),st6col44(1),st6col44(2),st5col44(4),st5col45(0));
fa1st6col44: FA port map(st6col44(3),st6col44(4),st6col44(5),st5col44(5),st5col45(1));
fa2st6col44: FA port map(st6col44(6),st6col44(7),st6col44(8),st5col44(6),st5col45(2));
fa3st6col44: FA port map(st6col44(9),st6col44(10),st6col44(11),st5col44(7),st5col45(3));
st5col44(8)<=st6col44(12);
fa0st6col45: FA port map(st6col45(0),st6col45(1),st6col45(2),st5col45(4),st5col46(0));
fa1st6col45: FA port map(st6col45(3),st6col45(4),st6col45(5),st5col45(5),st5col46(1));
fa2st6col45: FA port map(st6col45(6),st6col45(7),st6col45(8),st5col45(6),st5col46(2));
ha1st6col45: HA port map(st6col45(9),st6col45(10),st5col45(7),st5col46(3));
st5col45(8)<=st6col45(11);
fa0st6col46: FA port map(st6col46(0),st6col46(1),st6col46(2),st5col46(4),st5col47(0));
fa1st6col46: FA port map(st6col46(3),st6col46(4),st6col46(5),st5col46(5),st5col47(1));
fa2st6col46: FA port map(st6col46(6),st6col46(7),st6col46(8),st5col46(6),st5col47(2));
st5col46(7)<=st6col46(9);
st5col46(8)<=st6col46(10);
fa0st6col47: FA port map(st6col47(0),st6col47(1),st6col47(2),st5col47(3),st5col48(0));
fa1st6col47: FA port map(st6col47(3),st6col47(4),st6col47(5),st5col47(4),st5col48(1));
ha1st6col47: HA port map(st6col47(6),st6col47(7),st5col47(5),st5col48(2));
st5col47(6)<=st6col47(8);
st5col47(7)<=st6col47(9);
st5col47(8)<=st6col47(10);
fa0st6col48: FA port map(st6col48(0),st6col48(1),st6col48(2),st5col48(3),st5col49(0));
fa1st6col48: FA port map(st6col48(3),st6col48(4),st6col48(5),st5col48(4),st5col49(1));
st5col48(5)<=st6col48(6);
st5col48(6)<=st6col48(7);
st5col48(7)<=st6col48(8);
st5col48(8)<=st6col48(9);
fa0st6col49: FA port map(st6col49(0),st6col49(1),st6col49(2),st5col49(2),st5col50(0));
ha1st6col49: HA port map(st6col49(3),st6col49(4),st5col49(3),st5col50(1));
st5col49(4)<=st6col49(5);
st5col49(5)<=st6col49(6);
st5col49(6)<=st6col49(7);
st5col49(7)<=st6col49(8);
st5col49(8)<=st6col49(9);
fa0st6col50: FA port map(st6col50(0),st6col50(1),st6col50(2),st5col50(2),st5col51(0));
st5col50(3)<=st6col50(3);
st5col50(4)<=st6col50(4);
st5col50(5)<=st6col50(5);
st5col50(6)<=st6col50(6);
st5col50(7)<=st6col50(7);
st5col50(8)<=st6col50(8);
ha1st6col51: HA port map(st6col51(0),st6col51(1),st5col51(1),st5col52(0));
st5col51(2)<=st6col51(2);
st5col51(3)<=st6col51(3);
st5col51(4)<=st6col51(4);
st5col51(5)<=st6col51(5);
st5col51(6)<=st6col51(6);
st5col51(7)<=st6col51(7);
st5col51(8)<=st6col51(8);
st5col52(1)<=st6col52(0);
st5col52(2)<=st6col52(1);
st5col52(3)<=st6col52(2);
st5col52(4)<=st6col52(3);
st5col52(5)<=st6col52(4);
st5col52(6)<=st6col52(5);
st5col52(7)<=st6col52(6);
st5col52(8)<=st6col52(7);
st5col53(0)<=st6col53(0);
st5col53(1)<=st6col53(1);
st5col53(2)<=st6col53(2);
st5col53(3)<=st6col53(3);
st5col53(4)<=st6col53(4);
st5col53(5)<=st6col53(5);
st5col53(6)<=st6col53(6);
st5col53(7)<=st6col53(7);
st5col54(0)<=st6col54(0);
st5col54(1)<=st6col54(1);
st5col54(2)<=st6col54(2);
st5col54(3)<=st6col54(3);
st5col54(4)<=st6col54(4);
st5col54(5)<=st6col54(5);
st5col54(6)<=st6col54(6);
st5col55(0)<=st6col55(0);
st5col55(1)<=st6col55(1);
st5col55(2)<=st6col55(2);
st5col55(3)<=st6col55(3);
st5col55(4)<=st6col55(4);
st5col55(5)<=st6col55(5);
st5col55(6)<=st6col55(6);
st5col56(0)<=st6col56(0);
st5col56(1)<=st6col56(1);
st5col56(2)<=st6col56(2);
st5col56(3)<=st6col56(3);
st5col56(4)<=st6col56(4);
st5col56(5)<=st6col56(5);
st5col57(0)<=st6col57(0);
st5col57(1)<=st6col57(1);
st5col57(2)<=st6col57(2);
st5col57(3)<=st6col57(3);
st5col57(4)<=st6col57(4);
st5col57(5)<=st6col57(5);
st5col58(0)<=st6col58(0);
st5col58(1)<=st6col58(1);
st5col58(2)<=st6col58(2);
st5col58(3)<=st6col58(3);
st5col58(4)<=st6col58(4);
st5col59(0)<=st6col59(0);
st5col59(1)<=st6col59(1);
st5col59(2)<=st6col59(2);
st5col59(3)<=st6col59(3);
st5col59(4)<=st6col59(4);
st5col60(0)<=st6col60(0);
st5col60(1)<=st6col60(1);
st5col60(2)<=st6col60(2);
st5col60(3)<=st6col60(3);
st5col61(0)<=st6col61(0);
st5col61(1)<=st6col61(1);
st5col61(2)<=st6col61(2);
st5col61(3)<=st6col61(3);
st5col62(0)<=st6col62(0);
st5col62(1)<=st6col62(1);
st5col62(2)<=st6col62(2);
st5col63(0)<=st6col63(0);
st5col63(1)<=st6col63(1);
st5col63(2)<=st6col63(2);
st5col64(0)<=st6col64(0);
st5col64(1)<=st6col64(1);
st4col1(0)<=st5col1(0);
st4col1(1)<=st5col1(1);
st4col2(0)<=st5col2(0);
st4col3(0)<=st5col3(0);
st4col3(1)<=st5col3(1);
st4col3(2)<=st5col3(2);
st4col4(0)<=st5col4(0);
st4col4(1)<=st5col4(1);
st4col5(0)<=st5col5(0);
st4col5(1)<=st5col5(1);
st4col5(2)<=st5col5(2);
st4col5(3)<=st5col5(3);
st4col6(0)<=st5col6(0);
st4col6(1)<=st5col6(1);
st4col6(2)<=st5col6(2);
st4col7(0)<=st5col7(0);
st4col7(1)<=st5col7(1);
st4col7(2)<=st5col7(2);
st4col7(3)<=st5col7(3);
st4col7(4)<=st5col7(4);
st4col8(0)<=st5col8(0);
st4col8(1)<=st5col8(1);
st4col8(2)<=st5col8(2);
st4col8(3)<=st5col8(3);
st4col9(0)<=st5col9(0);
st4col9(1)<=st5col9(1);
st4col9(2)<=st5col9(2);
st4col9(3)<=st5col9(3);
st4col9(4)<=st5col9(4);
st4col9(5)<=st5col9(5);
st4col10(0)<=st5col10(0);
st4col10(1)<=st5col10(1);
st4col10(2)<=st5col10(2);
st4col10(3)<=st5col10(3);
st4col10(4)<=st5col10(4);
ha1st5col11: HA port map(st5col11(0),st5col11(1),st4col11(0),st4col12(0));
st4col11(1)<=st5col11(2);
st4col11(2)<=st5col11(3);
st4col11(3)<=st5col11(4);
st4col11(4)<=st5col11(5);
st4col11(5)<=st5col11(6);
ha1st5col12: HA port map(st5col12(0),st5col12(1),st4col12(1),st4col13(0));
st4col12(2)<=st5col12(2);
st4col12(3)<=st5col12(3);
st4col12(4)<=st5col12(4);
st4col12(5)<=st5col12(5);
fa0st5col13: FA port map(st5col13(0),st5col13(1),st5col13(2),st4col13(1),st4col14(0));
ha1st5col13: HA port map(st5col13(3),st5col13(4),st4col13(2),st4col14(1));
st4col13(3)<=st5col13(5);
st4col13(4)<=st5col13(6);
st4col13(5)<=st5col13(7);
fa0st5col14: FA port map(st5col14(0),st5col14(1),st5col14(2),st4col14(2),st4col15(0));
ha1st5col14: HA port map(st5col14(3),st5col14(4),st4col14(3),st4col15(1));
st4col14(4)<=st5col14(5);
st4col14(5)<=st5col14(6);
fa0st5col15: FA port map(st5col15(0),st5col15(1),st5col15(2),st4col15(2),st4col16(0));
fa1st5col15: FA port map(st5col15(3),st5col15(4),st5col15(5),st4col15(3),st4col16(1));
ha1st5col15: HA port map(st5col15(6),st5col15(7),st4col15(4),st4col16(2));
st4col15(5)<=st5col15(8);
fa0st5col16: FA port map(st5col16(0),st5col16(1),st5col16(2),st4col16(3),st4col17(0));
fa1st5col16: FA port map(st5col16(3),st5col16(4),st5col16(5),st4col16(4),st4col17(1));
ha1st5col16: HA port map(st5col16(6),st5col16(7),st4col16(5),st4col17(2));
fa0st5col17: FA port map(st5col17(0),st5col17(1),st5col17(2),st4col17(3),st4col18(0));
fa1st5col17: FA port map(st5col17(3),st5col17(4),st5col17(5),st4col17(4),st4col18(1));
fa2st5col17: FA port map(st5col17(6),st5col17(7),st5col17(8),st4col17(5),st4col18(2));
fa0st5col18: FA port map(st5col18(0),st5col18(1),st5col18(2),st4col18(3),st4col19(0));
fa1st5col18: FA port map(st5col18(3),st5col18(4),st5col18(5),st4col18(4),st4col19(1));
fa2st5col18: FA port map(st5col18(6),st5col18(7),st5col18(8),st4col18(5),st4col19(2));
fa0st5col19: FA port map(st5col19(0),st5col19(1),st5col19(2),st4col19(3),st4col20(0));
fa1st5col19: FA port map(st5col19(3),st5col19(4),st5col19(5),st4col19(4),st4col20(1));
fa2st5col19: FA port map(st5col19(6),st5col19(7),st5col19(8),st4col19(5),st4col20(2));
fa0st5col20: FA port map(st5col20(0),st5col20(1),st5col20(2),st4col20(3),st4col21(0));
fa1st5col20: FA port map(st5col20(3),st5col20(4),st5col20(5),st4col20(4),st4col21(1));
fa2st5col20: FA port map(st5col20(6),st5col20(7),st5col20(8),st4col20(5),st4col21(2));
fa0st5col21: FA port map(st5col21(0),st5col21(1),st5col21(2),st4col21(3),st4col22(0));
fa1st5col21: FA port map(st5col21(3),st5col21(4),st5col21(5),st4col21(4),st4col22(1));
fa2st5col21: FA port map(st5col21(6),st5col21(7),st5col21(8),st4col21(5),st4col22(2));
fa0st5col22: FA port map(st5col22(0),st5col22(1),st5col22(2),st4col22(3),st4col23(0));
fa1st5col22: FA port map(st5col22(3),st5col22(4),st5col22(5),st4col22(4),st4col23(1));
fa2st5col22: FA port map(st5col22(6),st5col22(7),st5col22(8),st4col22(5),st4col23(2));
fa0st5col23: FA port map(st5col23(0),st5col23(1),st5col23(2),st4col23(3),st4col24(0));
fa1st5col23: FA port map(st5col23(3),st5col23(4),st5col23(5),st4col23(4),st4col24(1));
fa2st5col23: FA port map(st5col23(6),st5col23(7),st5col23(8),st4col23(5),st4col24(2));
fa0st5col24: FA port map(st5col24(0),st5col24(1),st5col24(2),st4col24(3),st4col25(0));
fa1st5col24: FA port map(st5col24(3),st5col24(4),st5col24(5),st4col24(4),st4col25(1));
fa2st5col24: FA port map(st5col24(6),st5col24(7),st5col24(8),st4col24(5),st4col25(2));
fa0st5col25: FA port map(st5col25(0),st5col25(1),st5col25(2),st4col25(3),st4col26(0));
fa1st5col25: FA port map(st5col25(3),st5col25(4),st5col25(5),st4col25(4),st4col26(1));
fa2st5col25: FA port map(st5col25(6),st5col25(7),st5col25(8),st4col25(5),st4col26(2));
fa0st5col26: FA port map(st5col26(0),st5col26(1),st5col26(2),st4col26(3),st4col27(0));
fa1st5col26: FA port map(st5col26(3),st5col26(4),st5col26(5),st4col26(4),st4col27(1));
fa2st5col26: FA port map(st5col26(6),st5col26(7),st5col26(8),st4col26(5),st4col27(2));
fa0st5col27: FA port map(st5col27(0),st5col27(1),st5col27(2),st4col27(3),st4col28(0));
fa1st5col27: FA port map(st5col27(3),st5col27(4),st5col27(5),st4col27(4),st4col28(1));
fa2st5col27: FA port map(st5col27(6),st5col27(7),st5col27(8),st4col27(5),st4col28(2));
fa0st5col28: FA port map(st5col28(0),st5col28(1),st5col28(2),st4col28(3),st4col29(0));
fa1st5col28: FA port map(st5col28(3),st5col28(4),st5col28(5),st4col28(4),st4col29(1));
fa2st5col28: FA port map(st5col28(6),st5col28(7),st5col28(8),st4col28(5),st4col29(2));
fa0st5col29: FA port map(st5col29(0),st5col29(1),st5col29(2),st4col29(3),st4col30(0));
fa1st5col29: FA port map(st5col29(3),st5col29(4),st5col29(5),st4col29(4),st4col30(1));
fa2st5col29: FA port map(st5col29(6),st5col29(7),st5col29(8),st4col29(5),st4col30(2));
fa0st5col30: FA port map(st5col30(0),st5col30(1),st5col30(2),st4col30(3),st4col31(0));
fa1st5col30: FA port map(st5col30(3),st5col30(4),st5col30(5),st4col30(4),st4col31(1));
fa2st5col30: FA port map(st5col30(6),st5col30(7),st5col30(8),st4col30(5),st4col31(2));
fa0st5col31: FA port map(st5col31(0),st5col31(1),st5col31(2),st4col31(3),st4col32(0));
fa1st5col31: FA port map(st5col31(3),st5col31(4),st5col31(5),st4col31(4),st4col32(1));
fa2st5col31: FA port map(st5col31(6),st5col31(7),st5col31(8),st4col31(5),st4col32(2));
fa0st5col32: FA port map(st5col32(0),st5col32(1),st5col32(2),st4col32(3),st4col33(0));
fa1st5col32: FA port map(st5col32(3),st5col32(4),st5col32(5),st4col32(4),st4col33(1));
fa2st5col32: FA port map(st5col32(6),st5col32(7),st5col32(8),st4col32(5),st4col33(2));
fa0st5col33: FA port map(st5col33(0),st5col33(1),st5col33(2),st4col33(3),st4col34(0));
fa1st5col33: FA port map(st5col33(3),st5col33(4),st5col33(5),st4col33(4),st4col34(1));
fa2st5col33: FA port map(st5col33(6),st5col33(7),st5col33(8),st4col33(5),st4col34(2));
fa0st5col34: FA port map(st5col34(0),st5col34(1),st5col34(2),st4col34(3),st4col35(0));
fa1st5col34: FA port map(st5col34(3),st5col34(4),st5col34(5),st4col34(4),st4col35(1));
fa2st5col34: FA port map(st5col34(6),st5col34(7),st5col34(8),st4col34(5),st4col35(2));
fa0st5col35: FA port map(st5col35(0),st5col35(1),st5col35(2),st4col35(3),st4col36(0));
fa1st5col35: FA port map(st5col35(3),st5col35(4),st5col35(5),st4col35(4),st4col36(1));
fa2st5col35: FA port map(st5col35(6),st5col35(7),st5col35(8),st4col35(5),st4col36(2));
fa0st5col36: FA port map(st5col36(0),st5col36(1),st5col36(2),st4col36(3),st4col37(0));
fa1st5col36: FA port map(st5col36(3),st5col36(4),st5col36(5),st4col36(4),st4col37(1));
fa2st5col36: FA port map(st5col36(6),st5col36(7),st5col36(8),st4col36(5),st4col37(2));
fa0st5col37: FA port map(st5col37(0),st5col37(1),st5col37(2),st4col37(3),st4col38(0));
fa1st5col37: FA port map(st5col37(3),st5col37(4),st5col37(5),st4col37(4),st4col38(1));
fa2st5col37: FA port map(st5col37(6),st5col37(7),st5col37(8),st4col37(5),st4col38(2));
fa0st5col38: FA port map(st5col38(0),st5col38(1),st5col38(2),st4col38(3),st4col39(0));
fa1st5col38: FA port map(st5col38(3),st5col38(4),st5col38(5),st4col38(4),st4col39(1));
fa2st5col38: FA port map(st5col38(6),st5col38(7),st5col38(8),st4col38(5),st4col39(2));
fa0st5col39: FA port map(st5col39(0),st5col39(1),st5col39(2),st4col39(3),st4col40(0));
fa1st5col39: FA port map(st5col39(3),st5col39(4),st5col39(5),st4col39(4),st4col40(1));
fa2st5col39: FA port map(st5col39(6),st5col39(7),st5col39(8),st4col39(5),st4col40(2));
fa0st5col40: FA port map(st5col40(0),st5col40(1),st5col40(2),st4col40(3),st4col41(0));
fa1st5col40: FA port map(st5col40(3),st5col40(4),st5col40(5),st4col40(4),st4col41(1));
fa2st5col40: FA port map(st5col40(6),st5col40(7),st5col40(8),st4col40(5),st4col41(2));
fa0st5col41: FA port map(st5col41(0),st5col41(1),st5col41(2),st4col41(3),st4col42(0));
fa1st5col41: FA port map(st5col41(3),st5col41(4),st5col41(5),st4col41(4),st4col42(1));
fa2st5col41: FA port map(st5col41(6),st5col41(7),st5col41(8),st4col41(5),st4col42(2));
fa0st5col42: FA port map(st5col42(0),st5col42(1),st5col42(2),st4col42(3),st4col43(0));
fa1st5col42: FA port map(st5col42(3),st5col42(4),st5col42(5),st4col42(4),st4col43(1));
fa2st5col42: FA port map(st5col42(6),st5col42(7),st5col42(8),st4col42(5),st4col43(2));
fa0st5col43: FA port map(st5col43(0),st5col43(1),st5col43(2),st4col43(3),st4col44(0));
fa1st5col43: FA port map(st5col43(3),st5col43(4),st5col43(5),st4col43(4),st4col44(1));
fa2st5col43: FA port map(st5col43(6),st5col43(7),st5col43(8),st4col43(5),st4col44(2));
fa0st5col44: FA port map(st5col44(0),st5col44(1),st5col44(2),st4col44(3),st4col45(0));
fa1st5col44: FA port map(st5col44(3),st5col44(4),st5col44(5),st4col44(4),st4col45(1));
fa2st5col44: FA port map(st5col44(6),st5col44(7),st5col44(8),st4col44(5),st4col45(2));
fa0st5col45: FA port map(st5col45(0),st5col45(1),st5col45(2),st4col45(3),st4col46(0));
fa1st5col45: FA port map(st5col45(3),st5col45(4),st5col45(5),st4col45(4),st4col46(1));
fa2st5col45: FA port map(st5col45(6),st5col45(7),st5col45(8),st4col45(5),st4col46(2));
fa0st5col46: FA port map(st5col46(0),st5col46(1),st5col46(2),st4col46(3),st4col47(0));
fa1st5col46: FA port map(st5col46(3),st5col46(4),st5col46(5),st4col46(4),st4col47(1));
fa2st5col46: FA port map(st5col46(6),st5col46(7),st5col46(8),st4col46(5),st4col47(2));
fa0st5col47: FA port map(st5col47(0),st5col47(1),st5col47(2),st4col47(3),st4col48(0));
fa1st5col47: FA port map(st5col47(3),st5col47(4),st5col47(5),st4col47(4),st4col48(1));
fa2st5col47: FA port map(st5col47(6),st5col47(7),st5col47(8),st4col47(5),st4col48(2));
fa0st5col48: FA port map(st5col48(0),st5col48(1),st5col48(2),st4col48(3),st4col49(0));
fa1st5col48: FA port map(st5col48(3),st5col48(4),st5col48(5),st4col48(4),st4col49(1));
fa2st5col48: FA port map(st5col48(6),st5col48(7),st5col48(8),st4col48(5),st4col49(2));
fa0st5col49: FA port map(st5col49(0),st5col49(1),st5col49(2),st4col49(3),st4col50(0));
fa1st5col49: FA port map(st5col49(3),st5col49(4),st5col49(5),st4col49(4),st4col50(1));
fa2st5col49: FA port map(st5col49(6),st5col49(7),st5col49(8),st4col49(5),st4col50(2));
fa0st5col50: FA port map(st5col50(0),st5col50(1),st5col50(2),st4col50(3),st4col51(0));
fa1st5col50: FA port map(st5col50(3),st5col50(4),st5col50(5),st4col50(4),st4col51(1));
fa2st5col50: FA port map(st5col50(6),st5col50(7),st5col50(8),st4col50(5),st4col51(2));
fa0st5col51: FA port map(st5col51(0),st5col51(1),st5col51(2),st4col51(3),st4col52(0));
fa1st5col51: FA port map(st5col51(3),st5col51(4),st5col51(5),st4col51(4),st4col52(1));
fa2st5col51: FA port map(st5col51(6),st5col51(7),st5col51(8),st4col51(5),st4col52(2));
fa0st5col52: FA port map(st5col52(0),st5col52(1),st5col52(2),st4col52(3),st4col53(0));
fa1st5col52: FA port map(st5col52(3),st5col52(4),st5col52(5),st4col52(4),st4col53(1));
fa2st5col52: FA port map(st5col52(6),st5col52(7),st5col52(8),st4col52(5),st4col53(2));
fa0st5col53: FA port map(st5col53(0),st5col53(1),st5col53(2),st4col53(3),st4col54(0));
fa1st5col53: FA port map(st5col53(3),st5col53(4),st5col53(5),st4col53(4),st4col54(1));
ha1st5col53: HA port map(st5col53(6),st5col53(7),st4col53(5),st4col54(2));
fa0st5col54: FA port map(st5col54(0),st5col54(1),st5col54(2),st4col54(3),st4col55(0));
fa1st5col54: FA port map(st5col54(3),st5col54(4),st5col54(5),st4col54(4),st4col55(1));
st4col54(5)<=st5col54(6);
fa0st5col55: FA port map(st5col55(0),st5col55(1),st5col55(2),st4col55(2),st4col56(0));
ha1st5col55: HA port map(st5col55(3),st5col55(4),st4col55(3),st4col56(1));
st4col55(4)<=st5col55(5);
st4col55(5)<=st5col55(6);
fa0st5col56: FA port map(st5col56(0),st5col56(1),st5col56(2),st4col56(2),st4col57(0));
st4col56(3)<=st5col56(3);
st4col56(4)<=st5col56(4);
st4col56(5)<=st5col56(5);
ha1st5col57: HA port map(st5col57(0),st5col57(1),st4col57(1),st4col58(0));
st4col57(2)<=st5col57(2);
st4col57(3)<=st5col57(3);
st4col57(4)<=st5col57(4);
st4col57(5)<=st5col57(5);
st4col58(1)<=st5col58(0);
st4col58(2)<=st5col58(1);
st4col58(3)<=st5col58(2);
st4col58(4)<=st5col58(3);
st4col58(5)<=st5col58(4);
st4col59(0)<=st5col59(0);
st4col59(1)<=st5col59(1);
st4col59(2)<=st5col59(2);
st4col59(3)<=st5col59(3);
st4col59(4)<=st5col59(4);
st4col60(0)<=st5col60(0);
st4col60(1)<=st5col60(1);
st4col60(2)<=st5col60(2);
st4col60(3)<=st5col60(3);
st4col61(0)<=st5col61(0);
st4col61(1)<=st5col61(1);
st4col61(2)<=st5col61(2);
st4col61(3)<=st5col61(3);
st4col62(0)<=st5col62(0);
st4col62(1)<=st5col62(1);
st4col62(2)<=st5col62(2);
st4col63(0)<=st5col63(0);
st4col63(1)<=st5col63(1);
st4col63(2)<=st5col63(2);
st4col64(0)<=st5col64(0);
st4col64(1)<=st5col64(1);
st3col1(0)<=st4col1(0);
st3col1(1)<=st4col1(1);
st3col2(0)<=st4col2(0);
st3col3(0)<=st4col3(0);
st3col3(1)<=st4col3(1);
st3col3(2)<=st4col3(2);
st3col4(0)<=st4col4(0);
st3col4(1)<=st4col4(1);
st3col5(0)<=st4col5(0);
st3col5(1)<=st4col5(1);
st3col5(2)<=st4col5(2);
st3col5(3)<=st4col5(3);
st3col6(0)<=st4col6(0);
st3col6(1)<=st4col6(1);
st3col6(2)<=st4col6(2);
ha1st4col7: HA port map(st4col7(0),st4col7(1),st3col7(0),st3col8(0));
st3col7(1)<=st4col7(2);
st3col7(2)<=st4col7(3);
st3col7(3)<=st4col7(4);
ha1st4col8: HA port map(st4col8(0),st4col8(1),st3col8(1),st3col9(0));
st3col8(2)<=st4col8(2);
st3col8(3)<=st4col8(3);
fa0st4col9: FA port map(st4col9(0),st4col9(1),st4col9(2),st3col9(1),st3col10(0));
ha1st4col9: HA port map(st4col9(3),st4col9(4),st3col9(2),st3col10(1));
st3col9(3)<=st4col9(5);
fa0st4col10: FA port map(st4col10(0),st4col10(1),st4col10(2),st3col10(2),st3col11(0));
ha1st4col10: HA port map(st4col10(3),st4col10(4),st3col10(3),st3col11(1));
fa0st4col11: FA port map(st4col11(0),st4col11(1),st4col11(2),st3col11(2),st3col12(0));
fa1st4col11: FA port map(st4col11(3),st4col11(4),st4col11(5),st3col11(3),st3col12(1));
fa0st4col12: FA port map(st4col12(0),st4col12(1),st4col12(2),st3col12(2),st3col13(0));
fa1st4col12: FA port map(st4col12(3),st4col12(4),st4col12(5),st3col12(3),st3col13(1));
fa0st4col13: FA port map(st4col13(0),st4col13(1),st4col13(2),st3col13(2),st3col14(0));
fa1st4col13: FA port map(st4col13(3),st4col13(4),st4col13(5),st3col13(3),st3col14(1));
fa0st4col14: FA port map(st4col14(0),st4col14(1),st4col14(2),st3col14(2),st3col15(0));
fa1st4col14: FA port map(st4col14(3),st4col14(4),st4col14(5),st3col14(3),st3col15(1));
fa0st4col15: FA port map(st4col15(0),st4col15(1),st4col15(2),st3col15(2),st3col16(0));
fa1st4col15: FA port map(st4col15(3),st4col15(4),st4col15(5),st3col15(3),st3col16(1));
fa0st4col16: FA port map(st4col16(0),st4col16(1),st4col16(2),st3col16(2),st3col17(0));
fa1st4col16: FA port map(st4col16(3),st4col16(4),st4col16(5),st3col16(3),st3col17(1));
fa0st4col17: FA port map(st4col17(0),st4col17(1),st4col17(2),st3col17(2),st3col18(0));
fa1st4col17: FA port map(st4col17(3),st4col17(4),st4col17(5),st3col17(3),st3col18(1));
fa0st4col18: FA port map(st4col18(0),st4col18(1),st4col18(2),st3col18(2),st3col19(0));
fa1st4col18: FA port map(st4col18(3),st4col18(4),st4col18(5),st3col18(3),st3col19(1));
fa0st4col19: FA port map(st4col19(0),st4col19(1),st4col19(2),st3col19(2),st3col20(0));
fa1st4col19: FA port map(st4col19(3),st4col19(4),st4col19(5),st3col19(3),st3col20(1));
fa0st4col20: FA port map(st4col20(0),st4col20(1),st4col20(2),st3col20(2),st3col21(0));
fa1st4col20: FA port map(st4col20(3),st4col20(4),st4col20(5),st3col20(3),st3col21(1));
fa0st4col21: FA port map(st4col21(0),st4col21(1),st4col21(2),st3col21(2),st3col22(0));
fa1st4col21: FA port map(st4col21(3),st4col21(4),st4col21(5),st3col21(3),st3col22(1));
fa0st4col22: FA port map(st4col22(0),st4col22(1),st4col22(2),st3col22(2),st3col23(0));
fa1st4col22: FA port map(st4col22(3),st4col22(4),st4col22(5),st3col22(3),st3col23(1));
fa0st4col23: FA port map(st4col23(0),st4col23(1),st4col23(2),st3col23(2),st3col24(0));
fa1st4col23: FA port map(st4col23(3),st4col23(4),st4col23(5),st3col23(3),st3col24(1));
fa0st4col24: FA port map(st4col24(0),st4col24(1),st4col24(2),st3col24(2),st3col25(0));
fa1st4col24: FA port map(st4col24(3),st4col24(4),st4col24(5),st3col24(3),st3col25(1));
fa0st4col25: FA port map(st4col25(0),st4col25(1),st4col25(2),st3col25(2),st3col26(0));
fa1st4col25: FA port map(st4col25(3),st4col25(4),st4col25(5),st3col25(3),st3col26(1));
fa0st4col26: FA port map(st4col26(0),st4col26(1),st4col26(2),st3col26(2),st3col27(0));
fa1st4col26: FA port map(st4col26(3),st4col26(4),st4col26(5),st3col26(3),st3col27(1));
fa0st4col27: FA port map(st4col27(0),st4col27(1),st4col27(2),st3col27(2),st3col28(0));
fa1st4col27: FA port map(st4col27(3),st4col27(4),st4col27(5),st3col27(3),st3col28(1));
fa0st4col28: FA port map(st4col28(0),st4col28(1),st4col28(2),st3col28(2),st3col29(0));
fa1st4col28: FA port map(st4col28(3),st4col28(4),st4col28(5),st3col28(3),st3col29(1));
fa0st4col29: FA port map(st4col29(0),st4col29(1),st4col29(2),st3col29(2),st3col30(0));
fa1st4col29: FA port map(st4col29(3),st4col29(4),st4col29(5),st3col29(3),st3col30(1));
fa0st4col30: FA port map(st4col30(0),st4col30(1),st4col30(2),st3col30(2),st3col31(0));
fa1st4col30: FA port map(st4col30(3),st4col30(4),st4col30(5),st3col30(3),st3col31(1));
fa0st4col31: FA port map(st4col31(0),st4col31(1),st4col31(2),st3col31(2),st3col32(0));
fa1st4col31: FA port map(st4col31(3),st4col31(4),st4col31(5),st3col31(3),st3col32(1));
fa0st4col32: FA port map(st4col32(0),st4col32(1),st4col32(2),st3col32(2),st3col33(0));
fa1st4col32: FA port map(st4col32(3),st4col32(4),st4col32(5),st3col32(3),st3col33(1));
fa0st4col33: FA port map(st4col33(0),st4col33(1),st4col33(2),st3col33(2),st3col34(0));
fa1st4col33: FA port map(st4col33(3),st4col33(4),st4col33(5),st3col33(3),st3col34(1));
fa0st4col34: FA port map(st4col34(0),st4col34(1),st4col34(2),st3col34(2),st3col35(0));
fa1st4col34: FA port map(st4col34(3),st4col34(4),st4col34(5),st3col34(3),st3col35(1));
fa0st4col35: FA port map(st4col35(0),st4col35(1),st4col35(2),st3col35(2),st3col36(0));
fa1st4col35: FA port map(st4col35(3),st4col35(4),st4col35(5),st3col35(3),st3col36(1));
fa0st4col36: FA port map(st4col36(0),st4col36(1),st4col36(2),st3col36(2),st3col37(0));
fa1st4col36: FA port map(st4col36(3),st4col36(4),st4col36(5),st3col36(3),st3col37(1));
fa0st4col37: FA port map(st4col37(0),st4col37(1),st4col37(2),st3col37(2),st3col38(0));
fa1st4col37: FA port map(st4col37(3),st4col37(4),st4col37(5),st3col37(3),st3col38(1));
fa0st4col38: FA port map(st4col38(0),st4col38(1),st4col38(2),st3col38(2),st3col39(0));
fa1st4col38: FA port map(st4col38(3),st4col38(4),st4col38(5),st3col38(3),st3col39(1));
fa0st4col39: FA port map(st4col39(0),st4col39(1),st4col39(2),st3col39(2),st3col40(0));
fa1st4col39: FA port map(st4col39(3),st4col39(4),st4col39(5),st3col39(3),st3col40(1));
fa0st4col40: FA port map(st4col40(0),st4col40(1),st4col40(2),st3col40(2),st3col41(0));
fa1st4col40: FA port map(st4col40(3),st4col40(4),st4col40(5),st3col40(3),st3col41(1));
fa0st4col41: FA port map(st4col41(0),st4col41(1),st4col41(2),st3col41(2),st3col42(0));
fa1st4col41: FA port map(st4col41(3),st4col41(4),st4col41(5),st3col41(3),st3col42(1));
fa0st4col42: FA port map(st4col42(0),st4col42(1),st4col42(2),st3col42(2),st3col43(0));
fa1st4col42: FA port map(st4col42(3),st4col42(4),st4col42(5),st3col42(3),st3col43(1));
fa0st4col43: FA port map(st4col43(0),st4col43(1),st4col43(2),st3col43(2),st3col44(0));
fa1st4col43: FA port map(st4col43(3),st4col43(4),st4col43(5),st3col43(3),st3col44(1));
fa0st4col44: FA port map(st4col44(0),st4col44(1),st4col44(2),st3col44(2),st3col45(0));
fa1st4col44: FA port map(st4col44(3),st4col44(4),st4col44(5),st3col44(3),st3col45(1));
fa0st4col45: FA port map(st4col45(0),st4col45(1),st4col45(2),st3col45(2),st3col46(0));
fa1st4col45: FA port map(st4col45(3),st4col45(4),st4col45(5),st3col45(3),st3col46(1));
fa0st4col46: FA port map(st4col46(0),st4col46(1),st4col46(2),st3col46(2),st3col47(0));
fa1st4col46: FA port map(st4col46(3),st4col46(4),st4col46(5),st3col46(3),st3col47(1));
fa0st4col47: FA port map(st4col47(0),st4col47(1),st4col47(2),st3col47(2),st3col48(0));
fa1st4col47: FA port map(st4col47(3),st4col47(4),st4col47(5),st3col47(3),st3col48(1));
fa0st4col48: FA port map(st4col48(0),st4col48(1),st4col48(2),st3col48(2),st3col49(0));
fa1st4col48: FA port map(st4col48(3),st4col48(4),st4col48(5),st3col48(3),st3col49(1));
fa0st4col49: FA port map(st4col49(0),st4col49(1),st4col49(2),st3col49(2),st3col50(0));
fa1st4col49: FA port map(st4col49(3),st4col49(4),st4col49(5),st3col49(3),st3col50(1));
fa0st4col50: FA port map(st4col50(0),st4col50(1),st4col50(2),st3col50(2),st3col51(0));
fa1st4col50: FA port map(st4col50(3),st4col50(4),st4col50(5),st3col50(3),st3col51(1));
fa0st4col51: FA port map(st4col51(0),st4col51(1),st4col51(2),st3col51(2),st3col52(0));
fa1st4col51: FA port map(st4col51(3),st4col51(4),st4col51(5),st3col51(3),st3col52(1));
fa0st4col52: FA port map(st4col52(0),st4col52(1),st4col52(2),st3col52(2),st3col53(0));
fa1st4col52: FA port map(st4col52(3),st4col52(4),st4col52(5),st3col52(3),st3col53(1));
fa0st4col53: FA port map(st4col53(0),st4col53(1),st4col53(2),st3col53(2),st3col54(0));
fa1st4col53: FA port map(st4col53(3),st4col53(4),st4col53(5),st3col53(3),st3col54(1));
fa0st4col54: FA port map(st4col54(0),st4col54(1),st4col54(2),st3col54(2),st3col55(0));
fa1st4col54: FA port map(st4col54(3),st4col54(4),st4col54(5),st3col54(3),st3col55(1));
fa0st4col55: FA port map(st4col55(0),st4col55(1),st4col55(2),st3col55(2),st3col56(0));
fa1st4col55: FA port map(st4col55(3),st4col55(4),st4col55(5),st3col55(3),st3col56(1));
fa0st4col56: FA port map(st4col56(0),st4col56(1),st4col56(2),st3col56(2),st3col57(0));
fa1st4col56: FA port map(st4col56(3),st4col56(4),st4col56(5),st3col56(3),st3col57(1));
fa0st4col57: FA port map(st4col57(0),st4col57(1),st4col57(2),st3col57(2),st3col58(0));
fa1st4col57: FA port map(st4col57(3),st4col57(4),st4col57(5),st3col57(3),st3col58(1));
fa0st4col58: FA port map(st4col58(0),st4col58(1),st4col58(2),st3col58(2),st3col59(0));
fa1st4col58: FA port map(st4col58(3),st4col58(4),st4col58(5),st3col58(3),st3col59(1));
fa0st4col59: FA port map(st4col59(0),st4col59(1),st4col59(2),st3col59(2),st3col60(0));
ha1st4col59: HA port map(st4col59(3),st4col59(4),st3col59(3),st3col60(1));
fa0st4col60: FA port map(st4col60(0),st4col60(1),st4col60(2),st3col60(2),st3col61(0));
st3col60(3)<=st4col60(3);
ha1st4col61: HA port map(st4col61(0),st4col61(1),st3col61(1),st3col62(0));
st3col61(2)<=st4col61(2);
st3col61(3)<=st4col61(3);
st3col62(1)<=st4col62(0);
st3col62(2)<=st4col62(1);
st3col62(3)<=st4col62(2);
st3col63(0)<=st4col63(0);
st3col63(1)<=st4col63(1);
st3col63(2)<=st4col63(2);
st3col64(0)<=st4col64(0);
st3col64(1)<=st4col64(1);
st2col1(0)<=st3col1(0);
st2col1(1)<=st3col1(1);
st2col2(0)<=st3col2(0);
st2col3(0)<=st3col3(0);
st2col3(1)<=st3col3(1);
st2col3(2)<=st3col3(2);
st2col4(0)<=st3col4(0);
st2col4(1)<=st3col4(1);
ha1st3col5: HA port map(st3col5(0),st3col5(1),st2col5(0),st2col6(0));
st2col5(1)<=st3col5(2);
st2col5(2)<=st3col5(3);
ha1st3col6: HA port map(st3col6(0),st3col6(1),st2col6(1),st2col7(0));
st2col6(2)<=st3col6(2);
fa0st3col7: FA port map(st3col7(0),st3col7(1),st3col7(2),st2col7(1),st2col8(0));
st2col7(2)<=st3col7(3);
fa0st3col8: FA port map(st3col8(0),st3col8(1),st3col8(2),st2col8(1),st2col9(0));
st2col8(2)<=st3col8(3);
fa0st3col9: FA port map(st3col9(0),st3col9(1),st3col9(2),st2col9(1),st2col10(0));
st2col9(2)<=st3col9(3);
fa0st3col10: FA port map(st3col10(0),st3col10(1),st3col10(2),st2col10(1),st2col11(0));
st2col10(2)<=st3col10(3);
fa0st3col11: FA port map(st3col11(0),st3col11(1),st3col11(2),st2col11(1),st2col12(0));
st2col11(2)<=st3col11(3);
fa0st3col12: FA port map(st3col12(0),st3col12(1),st3col12(2),st2col12(1),st2col13(0));
st2col12(2)<=st3col12(3);
fa0st3col13: FA port map(st3col13(0),st3col13(1),st3col13(2),st2col13(1),st2col14(0));
st2col13(2)<=st3col13(3);
fa0st3col14: FA port map(st3col14(0),st3col14(1),st3col14(2),st2col14(1),st2col15(0));
st2col14(2)<=st3col14(3);
fa0st3col15: FA port map(st3col15(0),st3col15(1),st3col15(2),st2col15(1),st2col16(0));
st2col15(2)<=st3col15(3);
fa0st3col16: FA port map(st3col16(0),st3col16(1),st3col16(2),st2col16(1),st2col17(0));
st2col16(2)<=st3col16(3);
fa0st3col17: FA port map(st3col17(0),st3col17(1),st3col17(2),st2col17(1),st2col18(0));
st2col17(2)<=st3col17(3);
fa0st3col18: FA port map(st3col18(0),st3col18(1),st3col18(2),st2col18(1),st2col19(0));
st2col18(2)<=st3col18(3);
fa0st3col19: FA port map(st3col19(0),st3col19(1),st3col19(2),st2col19(1),st2col20(0));
st2col19(2)<=st3col19(3);
fa0st3col20: FA port map(st3col20(0),st3col20(1),st3col20(2),st2col20(1),st2col21(0));
st2col20(2)<=st3col20(3);
fa0st3col21: FA port map(st3col21(0),st3col21(1),st3col21(2),st2col21(1),st2col22(0));
st2col21(2)<=st3col21(3);
fa0st3col22: FA port map(st3col22(0),st3col22(1),st3col22(2),st2col22(1),st2col23(0));
st2col22(2)<=st3col22(3);
fa0st3col23: FA port map(st3col23(0),st3col23(1),st3col23(2),st2col23(1),st2col24(0));
st2col23(2)<=st3col23(3);
fa0st3col24: FA port map(st3col24(0),st3col24(1),st3col24(2),st2col24(1),st2col25(0));
st2col24(2)<=st3col24(3);
fa0st3col25: FA port map(st3col25(0),st3col25(1),st3col25(2),st2col25(1),st2col26(0));
st2col25(2)<=st3col25(3);
fa0st3col26: FA port map(st3col26(0),st3col26(1),st3col26(2),st2col26(1),st2col27(0));
st2col26(2)<=st3col26(3);
fa0st3col27: FA port map(st3col27(0),st3col27(1),st3col27(2),st2col27(1),st2col28(0));
st2col27(2)<=st3col27(3);
fa0st3col28: FA port map(st3col28(0),st3col28(1),st3col28(2),st2col28(1),st2col29(0));
st2col28(2)<=st3col28(3);
fa0st3col29: FA port map(st3col29(0),st3col29(1),st3col29(2),st2col29(1),st2col30(0));
st2col29(2)<=st3col29(3);
fa0st3col30: FA port map(st3col30(0),st3col30(1),st3col30(2),st2col30(1),st2col31(0));
st2col30(2)<=st3col30(3);
fa0st3col31: FA port map(st3col31(0),st3col31(1),st3col31(2),st2col31(1),st2col32(0));
st2col31(2)<=st3col31(3);
fa0st3col32: FA port map(st3col32(0),st3col32(1),st3col32(2),st2col32(1),st2col33(0));
st2col32(2)<=st3col32(3);
fa0st3col33: FA port map(st3col33(0),st3col33(1),st3col33(2),st2col33(1),st2col34(0));
st2col33(2)<=st3col33(3);
fa0st3col34: FA port map(st3col34(0),st3col34(1),st3col34(2),st2col34(1),st2col35(0));
st2col34(2)<=st3col34(3);
fa0st3col35: FA port map(st3col35(0),st3col35(1),st3col35(2),st2col35(1),st2col36(0));
st2col35(2)<=st3col35(3);
fa0st3col36: FA port map(st3col36(0),st3col36(1),st3col36(2),st2col36(1),st2col37(0));
st2col36(2)<=st3col36(3);
fa0st3col37: FA port map(st3col37(0),st3col37(1),st3col37(2),st2col37(1),st2col38(0));
st2col37(2)<=st3col37(3);
fa0st3col38: FA port map(st3col38(0),st3col38(1),st3col38(2),st2col38(1),st2col39(0));
st2col38(2)<=st3col38(3);
fa0st3col39: FA port map(st3col39(0),st3col39(1),st3col39(2),st2col39(1),st2col40(0));
st2col39(2)<=st3col39(3);
fa0st3col40: FA port map(st3col40(0),st3col40(1),st3col40(2),st2col40(1),st2col41(0));
st2col40(2)<=st3col40(3);
fa0st3col41: FA port map(st3col41(0),st3col41(1),st3col41(2),st2col41(1),st2col42(0));
st2col41(2)<=st3col41(3);
fa0st3col42: FA port map(st3col42(0),st3col42(1),st3col42(2),st2col42(1),st2col43(0));
st2col42(2)<=st3col42(3);
fa0st3col43: FA port map(st3col43(0),st3col43(1),st3col43(2),st2col43(1),st2col44(0));
st2col43(2)<=st3col43(3);
fa0st3col44: FA port map(st3col44(0),st3col44(1),st3col44(2),st2col44(1),st2col45(0));
st2col44(2)<=st3col44(3);
fa0st3col45: FA port map(st3col45(0),st3col45(1),st3col45(2),st2col45(1),st2col46(0));
st2col45(2)<=st3col45(3);
fa0st3col46: FA port map(st3col46(0),st3col46(1),st3col46(2),st2col46(1),st2col47(0));
st2col46(2)<=st3col46(3);
fa0st3col47: FA port map(st3col47(0),st3col47(1),st3col47(2),st2col47(1),st2col48(0));
st2col47(2)<=st3col47(3);
fa0st3col48: FA port map(st3col48(0),st3col48(1),st3col48(2),st2col48(1),st2col49(0));
st2col48(2)<=st3col48(3);
fa0st3col49: FA port map(st3col49(0),st3col49(1),st3col49(2),st2col49(1),st2col50(0));
st2col49(2)<=st3col49(3);
fa0st3col50: FA port map(st3col50(0),st3col50(1),st3col50(2),st2col50(1),st2col51(0));
st2col50(2)<=st3col50(3);
fa0st3col51: FA port map(st3col51(0),st3col51(1),st3col51(2),st2col51(1),st2col52(0));
st2col51(2)<=st3col51(3);
fa0st3col52: FA port map(st3col52(0),st3col52(1),st3col52(2),st2col52(1),st2col53(0));
st2col52(2)<=st3col52(3);
fa0st3col53: FA port map(st3col53(0),st3col53(1),st3col53(2),st2col53(1),st2col54(0));
st2col53(2)<=st3col53(3);
fa0st3col54: FA port map(st3col54(0),st3col54(1),st3col54(2),st2col54(1),st2col55(0));
st2col54(2)<=st3col54(3);
fa0st3col55: FA port map(st3col55(0),st3col55(1),st3col55(2),st2col55(1),st2col56(0));
st2col55(2)<=st3col55(3);
fa0st3col56: FA port map(st3col56(0),st3col56(1),st3col56(2),st2col56(1),st2col57(0));
st2col56(2)<=st3col56(3);
fa0st3col57: FA port map(st3col57(0),st3col57(1),st3col57(2),st2col57(1),st2col58(0));
st2col57(2)<=st3col57(3);
fa0st3col58: FA port map(st3col58(0),st3col58(1),st3col58(2),st2col58(1),st2col59(0));
st2col58(2)<=st3col58(3);
fa0st3col59: FA port map(st3col59(0),st3col59(1),st3col59(2),st2col59(1),st2col60(0));
st2col59(2)<=st3col59(3);
fa0st3col60: FA port map(st3col60(0),st3col60(1),st3col60(2),st2col60(1),st2col61(0));
st2col60(2)<=st3col60(3);
fa0st3col61: FA port map(st3col61(0),st3col61(1),st3col61(2),st2col61(1),st2col62(0));
st2col61(2)<=st3col61(3);
fa0st3col62: FA port map(st3col62(0),st3col62(1),st3col62(2),st2col62(1),st2col63(0));
st2col62(2)<=st3col62(3);
ha1st3col63: HA port map(st3col63(0),st3col63(1),st2col63(1),st2col64(0));
st2col63(2)<=st3col63(2);
st2col64(1)<=st3col64(0);
st2col64(2)<=st3col64(1);
st1col1(0)<=st2col1(0);
st1col1(1)<=st2col1(1);
st1col2(0)<=st2col2(0);
ha1st2col3: HA port map(st2col3(0),st2col3(1),st1col3(0),st1col4(0));
st1col3(1)<=st2col3(2);
ha1st2col4: HA port map(st2col4(0),st2col4(1),st1col4(1),st1col5(0));
fa0st2col5: FA port map(st2col5(0),st2col5(1),st2col5(2),st1col5(1),st1col6(0));
fa0st2col6: FA port map(st2col6(0),st2col6(1),st2col6(2),st1col6(1),st1col7(0));
fa0st2col7: FA port map(st2col7(0),st2col7(1),st2col7(2),st1col7(1),st1col8(0));
fa0st2col8: FA port map(st2col8(0),st2col8(1),st2col8(2),st1col8(1),st1col9(0));
fa0st2col9: FA port map(st2col9(0),st2col9(1),st2col9(2),st1col9(1),st1col10(0));
fa0st2col10: FA port map(st2col10(0),st2col10(1),st2col10(2),st1col10(1),st1col11(0));
fa0st2col11: FA port map(st2col11(0),st2col11(1),st2col11(2),st1col11(1),st1col12(0));
fa0st2col12: FA port map(st2col12(0),st2col12(1),st2col12(2),st1col12(1),st1col13(0));
fa0st2col13: FA port map(st2col13(0),st2col13(1),st2col13(2),st1col13(1),st1col14(0));
fa0st2col14: FA port map(st2col14(0),st2col14(1),st2col14(2),st1col14(1),st1col15(0));
fa0st2col15: FA port map(st2col15(0),st2col15(1),st2col15(2),st1col15(1),st1col16(0));
fa0st2col16: FA port map(st2col16(0),st2col16(1),st2col16(2),st1col16(1),st1col17(0));
fa0st2col17: FA port map(st2col17(0),st2col17(1),st2col17(2),st1col17(1),st1col18(0));
fa0st2col18: FA port map(st2col18(0),st2col18(1),st2col18(2),st1col18(1),st1col19(0));
fa0st2col19: FA port map(st2col19(0),st2col19(1),st2col19(2),st1col19(1),st1col20(0));
fa0st2col20: FA port map(st2col20(0),st2col20(1),st2col20(2),st1col20(1),st1col21(0));
fa0st2col21: FA port map(st2col21(0),st2col21(1),st2col21(2),st1col21(1),st1col22(0));
fa0st2col22: FA port map(st2col22(0),st2col22(1),st2col22(2),st1col22(1),st1col23(0));
fa0st2col23: FA port map(st2col23(0),st2col23(1),st2col23(2),st1col23(1),st1col24(0));
fa0st2col24: FA port map(st2col24(0),st2col24(1),st2col24(2),st1col24(1),st1col25(0));
fa0st2col25: FA port map(st2col25(0),st2col25(1),st2col25(2),st1col25(1),st1col26(0));
fa0st2col26: FA port map(st2col26(0),st2col26(1),st2col26(2),st1col26(1),st1col27(0));
fa0st2col27: FA port map(st2col27(0),st2col27(1),st2col27(2),st1col27(1),st1col28(0));
fa0st2col28: FA port map(st2col28(0),st2col28(1),st2col28(2),st1col28(1),st1col29(0));
fa0st2col29: FA port map(st2col29(0),st2col29(1),st2col29(2),st1col29(1),st1col30(0));
fa0st2col30: FA port map(st2col30(0),st2col30(1),st2col30(2),st1col30(1),st1col31(0));
fa0st2col31: FA port map(st2col31(0),st2col31(1),st2col31(2),st1col31(1),st1col32(0));
fa0st2col32: FA port map(st2col32(0),st2col32(1),st2col32(2),st1col32(1),st1col33(0));
fa0st2col33: FA port map(st2col33(0),st2col33(1),st2col33(2),st1col33(1),st1col34(0));
fa0st2col34: FA port map(st2col34(0),st2col34(1),st2col34(2),st1col34(1),st1col35(0));
fa0st2col35: FA port map(st2col35(0),st2col35(1),st2col35(2),st1col35(1),st1col36(0));
fa0st2col36: FA port map(st2col36(0),st2col36(1),st2col36(2),st1col36(1),st1col37(0));
fa0st2col37: FA port map(st2col37(0),st2col37(1),st2col37(2),st1col37(1),st1col38(0));
fa0st2col38: FA port map(st2col38(0),st2col38(1),st2col38(2),st1col38(1),st1col39(0));
fa0st2col39: FA port map(st2col39(0),st2col39(1),st2col39(2),st1col39(1),st1col40(0));
fa0st2col40: FA port map(st2col40(0),st2col40(1),st2col40(2),st1col40(1),st1col41(0));
fa0st2col41: FA port map(st2col41(0),st2col41(1),st2col41(2),st1col41(1),st1col42(0));
fa0st2col42: FA port map(st2col42(0),st2col42(1),st2col42(2),st1col42(1),st1col43(0));
fa0st2col43: FA port map(st2col43(0),st2col43(1),st2col43(2),st1col43(1),st1col44(0));
fa0st2col44: FA port map(st2col44(0),st2col44(1),st2col44(2),st1col44(1),st1col45(0));
fa0st2col45: FA port map(st2col45(0),st2col45(1),st2col45(2),st1col45(1),st1col46(0));
fa0st2col46: FA port map(st2col46(0),st2col46(1),st2col46(2),st1col46(1),st1col47(0));
fa0st2col47: FA port map(st2col47(0),st2col47(1),st2col47(2),st1col47(1),st1col48(0));
fa0st2col48: FA port map(st2col48(0),st2col48(1),st2col48(2),st1col48(1),st1col49(0));
fa0st2col49: FA port map(st2col49(0),st2col49(1),st2col49(2),st1col49(1),st1col50(0));
fa0st2col50: FA port map(st2col50(0),st2col50(1),st2col50(2),st1col50(1),st1col51(0));
fa0st2col51: FA port map(st2col51(0),st2col51(1),st2col51(2),st1col51(1),st1col52(0));
fa0st2col52: FA port map(st2col52(0),st2col52(1),st2col52(2),st1col52(1),st1col53(0));
fa0st2col53: FA port map(st2col53(0),st2col53(1),st2col53(2),st1col53(1),st1col54(0));
fa0st2col54: FA port map(st2col54(0),st2col54(1),st2col54(2),st1col54(1),st1col55(0));
fa0st2col55: FA port map(st2col55(0),st2col55(1),st2col55(2),st1col55(1),st1col56(0));
fa0st2col56: FA port map(st2col56(0),st2col56(1),st2col56(2),st1col56(1),st1col57(0));
fa0st2col57: FA port map(st2col57(0),st2col57(1),st2col57(2),st1col57(1),st1col58(0));
fa0st2col58: FA port map(st2col58(0),st2col58(1),st2col58(2),st1col58(1),st1col59(0));
fa0st2col59: FA port map(st2col59(0),st2col59(1),st2col59(2),st1col59(1),st1col60(0));
fa0st2col60: FA port map(st2col60(0),st2col60(1),st2col60(2),st1col60(1),st1col61(0));
fa0st2col61: FA port map(st2col61(0),st2col61(1),st2col61(2),st1col61(1),st1col62(0));
fa0st2col62: FA port map(st2col62(0),st2col62(1),st2col62(2),st1col62(1),st1col63(0));
fa0st2col63: FA port map(st2col63(0),st2col63(1),st2col63(2),st1col63(1),st1col64(0));
fa0st2col64: FA port map(st2col64(0),st2col64(1),st2col64(2),st1col64(1),open);
st7col1(0) <= pprod(0) (0);
st7col2(0) <= pprod(0) (1);
st7col3(0) <= pprod(0) (2);
st7col4(0) <= pprod(0) (3);
st7col5(0) <= pprod(0) (4);
st7col6(0) <= pprod(0) (5);
st7col7(0) <= pprod(0) (6);
st7col8(0) <= pprod(0) (7);
st7col9(0) <= pprod(0) (8);
st7col10(0) <= pprod(0) (9);
st7col11(0) <= pprod(0) (10);
st7col12(0) <= pprod(0) (11);
st7col13(0) <= pprod(0) (12);
st7col14(0) <= pprod(0) (13);
st7col15(0) <= pprod(0) (14);
st7col16(0) <= pprod(0) (15);
st7col17(0) <= pprod(0) (16);
st7col18(0) <= pprod(0) (17);
st7col19(0) <= pprod(0) (18);
st7col20(0) <= pprod(0) (19);
st7col21(0) <= pprod(0) (20);
st7col22(0) <= pprod(0) (21);
st7col23(0) <= pprod(0) (22);
st7col24(0) <= pprod(0) (23);
st7col25(0) <= pprod(0) (24);
st7col26(0) <= pprod(0) (25);
st7col27(0) <= pprod(0) (26);
st7col28(0) <= pprod(0) (27);
st7col29(0) <= pprod(0) (28);
st7col30(0) <= pprod(0) (29);
st7col31(0) <= pprod(0) (30);
st7col32(0) <= pprod(0) (31);
st7col33(0) <= pprod(0) (32);
st7col1(1) <= S(0);
st7col34(0) <= S(0);
st7col35(0) <= S(0);
st7col36(0) <= not S(0);
st7col3(1) <= pprod(1) (0);
st7col4(1) <= pprod(1) (1);
st7col5(1) <= pprod(1) (2);
st7col6(1) <= pprod(1) (3);
st7col7(1) <= pprod(1) (4);
st7col8(1) <= pprod(1) (5);
st7col9(1) <= pprod(1) (6);
st7col10(1) <= pprod(1) (7);
st7col11(1) <= pprod(1) (8);
st7col12(1) <= pprod(1) (9);
st7col13(1) <= pprod(1) (10);
st7col14(1) <= pprod(1) (11);
st7col15(1) <= pprod(1) (12);
st7col16(1) <= pprod(1) (13);
st7col17(1) <= pprod(1) (14);
st7col18(1) <= pprod(1) (15);
st7col19(1) <= pprod(1) (16);
st7col20(1) <= pprod(1) (17);
st7col21(1) <= pprod(1) (18);
st7col22(1) <= pprod(1) (19);
st7col23(1) <= pprod(1) (20);
st7col24(1) <= pprod(1) (21);
st7col25(1) <= pprod(1) (22);
st7col26(1) <= pprod(1) (23);
st7col27(1) <= pprod(1) (24);
st7col28(1) <= pprod(1) (25);
st7col29(1) <= pprod(1) (26);
st7col30(1) <= pprod(1) (27);
st7col31(1) <= pprod(1) (28);
st7col32(1) <= pprod(1) (29);
st7col33(1) <= pprod(1) (30);
st7col34(1) <= pprod(1) (31);
st7col35(1) <= pprod(1) (32);
st7col3(2) <= S(1);
st7col36(1) <= not S(1);
st7col37(0) <= '1';
st7col5(2) <= pprod(2) (0);
st7col6(2) <= pprod(2) (1);
st7col7(2) <= pprod(2) (2);
st7col8(2) <= pprod(2) (3);
st7col9(2) <= pprod(2) (4);
st7col10(2) <= pprod(2) (5);
st7col11(2) <= pprod(2) (6);
st7col12(2) <= pprod(2) (7);
st7col13(2) <= pprod(2) (8);
st7col14(2) <= pprod(2) (9);
st7col15(2) <= pprod(2) (10);
st7col16(2) <= pprod(2) (11);
st7col17(2) <= pprod(2) (12);
st7col18(2) <= pprod(2) (13);
st7col19(2) <= pprod(2) (14);
st7col20(2) <= pprod(2) (15);
st7col21(2) <= pprod(2) (16);
st7col22(2) <= pprod(2) (17);
st7col23(2) <= pprod(2) (18);
st7col24(2) <= pprod(2) (19);
st7col25(2) <= pprod(2) (20);
st7col26(2) <= pprod(2) (21);
st7col27(2) <= pprod(2) (22);
st7col28(2) <= pprod(2) (23);
st7col29(2) <= pprod(2) (24);
st7col30(2) <= pprod(2) (25);
st7col31(2) <= pprod(2) (26);
st7col32(2) <= pprod(2) (27);
st7col33(2) <= pprod(2) (28);
st7col34(2) <= pprod(2) (29);
st7col35(2) <= pprod(2) (30);
st7col36(2) <= pprod(2) (31);
st7col37(1) <= pprod(2) (32);
st7col5(3) <= S(2);
st7col38(0) <= not S(2);
st7col39(0) <= '1';
st7col7(3) <= pprod(3) (0);
st7col8(3) <= pprod(3) (1);
st7col9(3) <= pprod(3) (2);
st7col10(3) <= pprod(3) (3);
st7col11(3) <= pprod(3) (4);
st7col12(3) <= pprod(3) (5);
st7col13(3) <= pprod(3) (6);
st7col14(3) <= pprod(3) (7);
st7col15(3) <= pprod(3) (8);
st7col16(3) <= pprod(3) (9);
st7col17(3) <= pprod(3) (10);
st7col18(3) <= pprod(3) (11);
st7col19(3) <= pprod(3) (12);
st7col20(3) <= pprod(3) (13);
st7col21(3) <= pprod(3) (14);
st7col22(3) <= pprod(3) (15);
st7col23(3) <= pprod(3) (16);
st7col24(3) <= pprod(3) (17);
st7col25(3) <= pprod(3) (18);
st7col26(3) <= pprod(3) (19);
st7col27(3) <= pprod(3) (20);
st7col28(3) <= pprod(3) (21);
st7col29(3) <= pprod(3) (22);
st7col30(3) <= pprod(3) (23);
st7col31(3) <= pprod(3) (24);
st7col32(3) <= pprod(3) (25);
st7col33(3) <= pprod(3) (26);
st7col34(3) <= pprod(3) (27);
st7col35(3) <= pprod(3) (28);
st7col36(3) <= pprod(3) (29);
st7col37(2) <= pprod(3) (30);
st7col38(1) <= pprod(3) (31);
st7col39(1) <= pprod(3) (32);
st7col7(4) <= S(3);
st7col40(0) <= not S(3);
st7col41(0) <= '1';
st7col9(4) <= pprod(4) (0);
st7col10(4) <= pprod(4) (1);
st7col11(4) <= pprod(4) (2);
st7col12(4) <= pprod(4) (3);
st7col13(4) <= pprod(4) (4);
st7col14(4) <= pprod(4) (5);
st7col15(4) <= pprod(4) (6);
st7col16(4) <= pprod(4) (7);
st7col17(4) <= pprod(4) (8);
st7col18(4) <= pprod(4) (9);
st7col19(4) <= pprod(4) (10);
st7col20(4) <= pprod(4) (11);
st7col21(4) <= pprod(4) (12);
st7col22(4) <= pprod(4) (13);
st7col23(4) <= pprod(4) (14);
st7col24(4) <= pprod(4) (15);
st7col25(4) <= pprod(4) (16);
st7col26(4) <= pprod(4) (17);
st7col27(4) <= pprod(4) (18);
st7col28(4) <= pprod(4) (19);
st7col29(4) <= pprod(4) (20);
st7col30(4) <= pprod(4) (21);
st7col31(4) <= pprod(4) (22);
st7col32(4) <= pprod(4) (23);
st7col33(4) <= pprod(4) (24);
st7col34(4) <= pprod(4) (25);
st7col35(4) <= pprod(4) (26);
st7col36(4) <= pprod(4) (27);
st7col37(3) <= pprod(4) (28);
st7col38(2) <= pprod(4) (29);
st7col39(2) <= pprod(4) (30);
st7col40(1) <= pprod(4) (31);
st7col41(1) <= pprod(4) (32);
st7col9(5) <= S(4);
st7col42(0) <= not S(4);
st7col43(0) <= '1';
st7col11(5) <= pprod(5) (0);
st7col12(5) <= pprod(5) (1);
st7col13(5) <= pprod(5) (2);
st7col14(5) <= pprod(5) (3);
st7col15(5) <= pprod(5) (4);
st7col16(5) <= pprod(5) (5);
st7col17(5) <= pprod(5) (6);
st7col18(5) <= pprod(5) (7);
st7col19(5) <= pprod(5) (8);
st7col20(5) <= pprod(5) (9);
st7col21(5) <= pprod(5) (10);
st7col22(5) <= pprod(5) (11);
st7col23(5) <= pprod(5) (12);
st7col24(5) <= pprod(5) (13);
st7col25(5) <= pprod(5) (14);
st7col26(5) <= pprod(5) (15);
st7col27(5) <= pprod(5) (16);
st7col28(5) <= pprod(5) (17);
st7col29(5) <= pprod(5) (18);
st7col30(5) <= pprod(5) (19);
st7col31(5) <= pprod(5) (20);
st7col32(5) <= pprod(5) (21);
st7col33(5) <= pprod(5) (22);
st7col34(5) <= pprod(5) (23);
st7col35(5) <= pprod(5) (24);
st7col36(5) <= pprod(5) (25);
st7col37(4) <= pprod(5) (26);
st7col38(3) <= pprod(5) (27);
st7col39(3) <= pprod(5) (28);
st7col40(2) <= pprod(5) (29);
st7col41(2) <= pprod(5) (30);
st7col42(1) <= pprod(5) (31);
st7col43(1) <= pprod(5) (32);
st7col11(6) <= S(5);
st7col44(0) <= not S(5);
st7col45(0) <= '1';
st7col13(6) <= pprod(6) (0);
st7col14(6) <= pprod(6) (1);
st7col15(6) <= pprod(6) (2);
st7col16(6) <= pprod(6) (3);
st7col17(6) <= pprod(6) (4);
st7col18(6) <= pprod(6) (5);
st7col19(6) <= pprod(6) (6);
st7col20(6) <= pprod(6) (7);
st7col21(6) <= pprod(6) (8);
st7col22(6) <= pprod(6) (9);
st7col23(6) <= pprod(6) (10);
st7col24(6) <= pprod(6) (11);
st7col25(6) <= pprod(6) (12);
st7col26(6) <= pprod(6) (13);
st7col27(6) <= pprod(6) (14);
st7col28(6) <= pprod(6) (15);
st7col29(6) <= pprod(6) (16);
st7col30(6) <= pprod(6) (17);
st7col31(6) <= pprod(6) (18);
st7col32(6) <= pprod(6) (19);
st7col33(6) <= pprod(6) (20);
st7col34(6) <= pprod(6) (21);
st7col35(6) <= pprod(6) (22);
st7col36(6) <= pprod(6) (23);
st7col37(5) <= pprod(6) (24);
st7col38(4) <= pprod(6) (25);
st7col39(4) <= pprod(6) (26);
st7col40(3) <= pprod(6) (27);
st7col41(3) <= pprod(6) (28);
st7col42(2) <= pprod(6) (29);
st7col43(2) <= pprod(6) (30);
st7col44(1) <= pprod(6) (31);
st7col45(1) <= pprod(6) (32);
st7col13(7) <= S(6);
st7col46(0) <= not S(6);
st7col47(0) <= '1';
st7col15(7) <= pprod(7) (0);
st7col16(7) <= pprod(7) (1);
st7col17(7) <= pprod(7) (2);
st7col18(7) <= pprod(7) (3);
st7col19(7) <= pprod(7) (4);
st7col20(7) <= pprod(7) (5);
st7col21(7) <= pprod(7) (6);
st7col22(7) <= pprod(7) (7);
st7col23(7) <= pprod(7) (8);
st7col24(7) <= pprod(7) (9);
st7col25(7) <= pprod(7) (10);
st7col26(7) <= pprod(7) (11);
st7col27(7) <= pprod(7) (12);
st7col28(7) <= pprod(7) (13);
st7col29(7) <= pprod(7) (14);
st7col30(7) <= pprod(7) (15);
st7col31(7) <= pprod(7) (16);
st7col32(7) <= pprod(7) (17);
st7col33(7) <= pprod(7) (18);
st7col34(7) <= pprod(7) (19);
st7col35(7) <= pprod(7) (20);
st7col36(7) <= pprod(7) (21);
st7col37(6) <= pprod(7) (22);
st7col38(5) <= pprod(7) (23);
st7col39(5) <= pprod(7) (24);
st7col40(4) <= pprod(7) (25);
st7col41(4) <= pprod(7) (26);
st7col42(3) <= pprod(7) (27);
st7col43(3) <= pprod(7) (28);
st7col44(2) <= pprod(7) (29);
st7col45(2) <= pprod(7) (30);
st7col46(1) <= pprod(7) (31);
st7col47(1) <= pprod(7) (32);
st7col15(8) <= S(7);
st7col48(0) <= not S(7);
st7col49(0) <= '1';
st7col17(8) <= pprod(8) (0);
st7col18(8) <= pprod(8) (1);
st7col19(8) <= pprod(8) (2);
st7col20(8) <= pprod(8) (3);
st7col21(8) <= pprod(8) (4);
st7col22(8) <= pprod(8) (5);
st7col23(8) <= pprod(8) (6);
st7col24(8) <= pprod(8) (7);
st7col25(8) <= pprod(8) (8);
st7col26(8) <= pprod(8) (9);
st7col27(8) <= pprod(8) (10);
st7col28(8) <= pprod(8) (11);
st7col29(8) <= pprod(8) (12);
st7col30(8) <= pprod(8) (13);
st7col31(8) <= pprod(8) (14);
st7col32(8) <= pprod(8) (15);
st7col33(8) <= pprod(8) (16);
st7col34(8) <= pprod(8) (17);
st7col35(8) <= pprod(8) (18);
st7col36(8) <= pprod(8) (19);
st7col37(7) <= pprod(8) (20);
st7col38(6) <= pprod(8) (21);
st7col39(6) <= pprod(8) (22);
st7col40(5) <= pprod(8) (23);
st7col41(5) <= pprod(8) (24);
st7col42(4) <= pprod(8) (25);
st7col43(4) <= pprod(8) (26);
st7col44(3) <= pprod(8) (27);
st7col45(3) <= pprod(8) (28);
st7col46(2) <= pprod(8) (29);
st7col47(2) <= pprod(8) (30);
st7col48(1) <= pprod(8) (31);
st7col49(1) <= pprod(8) (32);
st7col17(9) <= S(8);
st7col50(0) <= not S(8);
st7col51(0) <= '1';
st7col19(9) <= pprod(9) (0);
st7col20(9) <= pprod(9) (1);
st7col21(9) <= pprod(9) (2);
st7col22(9) <= pprod(9) (3);
st7col23(9) <= pprod(9) (4);
st7col24(9) <= pprod(9) (5);
st7col25(9) <= pprod(9) (6);
st7col26(9) <= pprod(9) (7);
st7col27(9) <= pprod(9) (8);
st7col28(9) <= pprod(9) (9);
st7col29(9) <= pprod(9) (10);
st7col30(9) <= pprod(9) (11);
st7col31(9) <= pprod(9) (12);
st7col32(9) <= pprod(9) (13);
st7col33(9) <= pprod(9) (14);
st7col34(9) <= pprod(9) (15);
st7col35(9) <= pprod(9) (16);
st7col36(9) <= pprod(9) (17);
st7col37(8) <= pprod(9) (18);
st7col38(7) <= pprod(9) (19);
st7col39(7) <= pprod(9) (20);
st7col40(6) <= pprod(9) (21);
st7col41(6) <= pprod(9) (22);
st7col42(5) <= pprod(9) (23);
st7col43(5) <= pprod(9) (24);
st7col44(4) <= pprod(9) (25);
st7col45(4) <= pprod(9) (26);
st7col46(3) <= pprod(9) (27);
st7col47(3) <= pprod(9) (28);
st7col48(2) <= pprod(9) (29);
st7col49(2) <= pprod(9) (30);
st7col50(1) <= pprod(9) (31);
st7col51(1) <= pprod(9) (32);
st7col19(10) <= S(9);
st7col52(0) <= not S(9);
st7col53(0) <= '1';
st7col21(10) <= pprod(10) (0);
st7col22(10) <= pprod(10) (1);
st7col23(10) <= pprod(10) (2);
st7col24(10) <= pprod(10) (3);
st7col25(10) <= pprod(10) (4);
st7col26(10) <= pprod(10) (5);
st7col27(10) <= pprod(10) (6);
st7col28(10) <= pprod(10) (7);
st7col29(10) <= pprod(10) (8);
st7col30(10) <= pprod(10) (9);
st7col31(10) <= pprod(10) (10);
st7col32(10) <= pprod(10) (11);
st7col33(10) <= pprod(10) (12);
st7col34(10) <= pprod(10) (13);
st7col35(10) <= pprod(10) (14);
st7col36(10) <= pprod(10) (15);
st7col37(9) <= pprod(10) (16);
st7col38(8) <= pprod(10) (17);
st7col39(8) <= pprod(10) (18);
st7col40(7) <= pprod(10) (19);
st7col41(7) <= pprod(10) (20);
st7col42(6) <= pprod(10) (21);
st7col43(6) <= pprod(10) (22);
st7col44(5) <= pprod(10) (23);
st7col45(5) <= pprod(10) (24);
st7col46(4) <= pprod(10) (25);
st7col47(4) <= pprod(10) (26);
st7col48(3) <= pprod(10) (27);
st7col49(3) <= pprod(10) (28);
st7col50(2) <= pprod(10) (29);
st7col51(2) <= pprod(10) (30);
st7col52(1) <= pprod(10) (31);
st7col53(1) <= pprod(10) (32);
st7col21(11) <= S(10);
st7col54(0) <= not S(10);
st7col55(0) <= '1';
st7col23(11) <= pprod(11) (0);
st7col24(11) <= pprod(11) (1);
st7col25(11) <= pprod(11) (2);
st7col26(11) <= pprod(11) (3);
st7col27(11) <= pprod(11) (4);
st7col28(11) <= pprod(11) (5);
st7col29(11) <= pprod(11) (6);
st7col30(11) <= pprod(11) (7);
st7col31(11) <= pprod(11) (8);
st7col32(11) <= pprod(11) (9);
st7col33(11) <= pprod(11) (10);
st7col34(11) <= pprod(11) (11);
st7col35(11) <= pprod(11) (12);
st7col36(11) <= pprod(11) (13);
st7col37(10) <= pprod(11) (14);
st7col38(9) <= pprod(11) (15);
st7col39(9) <= pprod(11) (16);
st7col40(8) <= pprod(11) (17);
st7col41(8) <= pprod(11) (18);
st7col42(7) <= pprod(11) (19);
st7col43(7) <= pprod(11) (20);
st7col44(6) <= pprod(11) (21);
st7col45(6) <= pprod(11) (22);
st7col46(5) <= pprod(11) (23);
st7col47(5) <= pprod(11) (24);
st7col48(4) <= pprod(11) (25);
st7col49(4) <= pprod(11) (26);
st7col50(3) <= pprod(11) (27);
st7col51(3) <= pprod(11) (28);
st7col52(2) <= pprod(11) (29);
st7col53(2) <= pprod(11) (30);
st7col54(1) <= pprod(11) (31);
st7col55(1) <= pprod(11) (32);
st7col23(12) <= S(11);
st7col56(0) <= not S(11);
st7col57(0) <= '1';
st7col25(12) <= pprod(12) (0);
st7col26(12) <= pprod(12) (1);
st7col27(12) <= pprod(12) (2);
st7col28(12) <= pprod(12) (3);
st7col29(12) <= pprod(12) (4);
st7col30(12) <= pprod(12) (5);
st7col31(12) <= pprod(12) (6);
st7col32(12) <= pprod(12) (7);
st7col33(12) <= pprod(12) (8);
st7col34(12) <= pprod(12) (9);
st7col35(12) <= pprod(12) (10);
st7col36(12) <= pprod(12) (11);
st7col37(11) <= pprod(12) (12);
st7col38(10) <= pprod(12) (13);
st7col39(10) <= pprod(12) (14);
st7col40(9) <= pprod(12) (15);
st7col41(9) <= pprod(12) (16);
st7col42(8) <= pprod(12) (17);
st7col43(8) <= pprod(12) (18);
st7col44(7) <= pprod(12) (19);
st7col45(7) <= pprod(12) (20);
st7col46(6) <= pprod(12) (21);
st7col47(6) <= pprod(12) (22);
st7col48(5) <= pprod(12) (23);
st7col49(5) <= pprod(12) (24);
st7col50(4) <= pprod(12) (25);
st7col51(4) <= pprod(12) (26);
st7col52(3) <= pprod(12) (27);
st7col53(3) <= pprod(12) (28);
st7col54(2) <= pprod(12) (29);
st7col55(2) <= pprod(12) (30);
st7col56(1) <= pprod(12) (31);
st7col57(1) <= pprod(12) (32);
st7col25(13) <= S(12);
st7col58(0) <= not S(12);
st7col59(0) <= '1';
st7col27(13) <= pprod(13) (0);
st7col28(13) <= pprod(13) (1);
st7col29(13) <= pprod(13) (2);
st7col30(13) <= pprod(13) (3);
st7col31(13) <= pprod(13) (4);
st7col32(13) <= pprod(13) (5);
st7col33(13) <= pprod(13) (6);
st7col34(13) <= pprod(13) (7);
st7col35(13) <= pprod(13) (8);
st7col36(13) <= pprod(13) (9);
st7col37(12) <= pprod(13) (10);
st7col38(11) <= pprod(13) (11);
st7col39(11) <= pprod(13) (12);
st7col40(10) <= pprod(13) (13);
st7col41(10) <= pprod(13) (14);
st7col42(9) <= pprod(13) (15);
st7col43(9) <= pprod(13) (16);
st7col44(8) <= pprod(13) (17);
st7col45(8) <= pprod(13) (18);
st7col46(7) <= pprod(13) (19);
st7col47(7) <= pprod(13) (20);
st7col48(6) <= pprod(13) (21);
st7col49(6) <= pprod(13) (22);
st7col50(5) <= pprod(13) (23);
st7col51(5) <= pprod(13) (24);
st7col52(4) <= pprod(13) (25);
st7col53(4) <= pprod(13) (26);
st7col54(3) <= pprod(13) (27);
st7col55(3) <= pprod(13) (28);
st7col56(2) <= pprod(13) (29);
st7col57(2) <= pprod(13) (30);
st7col58(1) <= pprod(13) (31);
st7col59(1) <= pprod(13) (32);
st7col27(14) <= S(13);
st7col60(0) <= not S(13);
st7col61(0) <= '1';
st7col29(14) <= pprod(14) (0);
st7col30(14) <= pprod(14) (1);
st7col31(14) <= pprod(14) (2);
st7col32(14) <= pprod(14) (3);
st7col33(14) <= pprod(14) (4);
st7col34(14) <= pprod(14) (5);
st7col35(14) <= pprod(14) (6);
st7col36(14) <= pprod(14) (7);
st7col37(13) <= pprod(14) (8);
st7col38(12) <= pprod(14) (9);
st7col39(12) <= pprod(14) (10);
st7col40(11) <= pprod(14) (11);
st7col41(11) <= pprod(14) (12);
st7col42(10) <= pprod(14) (13);
st7col43(10) <= pprod(14) (14);
st7col44(9) <= pprod(14) (15);
st7col45(9) <= pprod(14) (16);
st7col46(8) <= pprod(14) (17);
st7col47(8) <= pprod(14) (18);
st7col48(7) <= pprod(14) (19);
st7col49(7) <= pprod(14) (20);
st7col50(6) <= pprod(14) (21);
st7col51(6) <= pprod(14) (22);
st7col52(5) <= pprod(14) (23);
st7col53(5) <= pprod(14) (24);
st7col54(4) <= pprod(14) (25);
st7col55(4) <= pprod(14) (26);
st7col56(3) <= pprod(14) (27);
st7col57(3) <= pprod(14) (28);
st7col58(2) <= pprod(14) (29);
st7col59(2) <= pprod(14) (30);
st7col60(1) <= pprod(14) (31);
st7col61(1) <= pprod(14) (32);
st7col29(15) <= S(14);
st7col62(0) <= not S(14);
st7col63(0) <= '1';
st7col31(15) <= pprod(15) (0);
st7col32(15) <= pprod(15) (1);
st7col33(15) <= pprod(15) (2);
st7col34(15) <= pprod(15) (3);
st7col35(15) <= pprod(15) (4);
st7col36(15) <= pprod(15) (5);
st7col37(14) <= pprod(15) (6);
st7col38(13) <= pprod(15) (7);
st7col39(13) <= pprod(15) (8);
st7col40(12) <= pprod(15) (9);
st7col41(12) <= pprod(15) (10);
st7col42(11) <= pprod(15) (11);
st7col43(11) <= pprod(15) (12);
st7col44(10) <= pprod(15) (13);
st7col45(10) <= pprod(15) (14);
st7col46(9) <= pprod(15) (15);
st7col47(9) <= pprod(15) (16);
st7col48(8) <= pprod(15) (17);
st7col49(8) <= pprod(15) (18);
st7col50(7) <= pprod(15) (19);
st7col51(7) <= pprod(15) (20);
st7col52(6) <= pprod(15) (21);
st7col53(6) <= pprod(15) (22);
st7col54(5) <= pprod(15) (23);
st7col55(5) <= pprod(15) (24);
st7col56(4) <= pprod(15) (25);
st7col57(4) <= pprod(15) (26);
st7col58(3) <= pprod(15) (27);
st7col59(3) <= pprod(15) (28);
st7col60(2) <= pprod(15) (29);
st7col61(2) <= pprod(15) (30);
st7col62(1) <= pprod(15) (31);
st7col63(1) <= pprod(15) (32);
st7col31(16) <= S(15);
st7col64(0) <= not S(15);
st7col33(16) <= pprod(16) (0);
st7col34(16) <= pprod(16) (1);
st7col35(16) <= pprod(16) (2);
st7col36(16) <= pprod(16) (3);
st7col37(15) <= pprod(16) (4);
st7col38(14) <= pprod(16) (5);
st7col39(14) <= pprod(16) (6);
st7col40(13) <= pprod(16) (7);
st7col41(13) <= pprod(16) (8);
st7col42(12) <= pprod(16) (9);
st7col43(12) <= pprod(16) (10);
st7col44(11) <= pprod(16) (11);
st7col45(11) <= pprod(16) (12);
st7col46(10) <= pprod(16) (13);
st7col47(10) <= pprod(16) (14);
st7col48(9) <= pprod(16) (15);
st7col49(9) <= pprod(16) (16);
st7col50(8) <= pprod(16) (17);
st7col51(8) <= pprod(16) (18);
st7col52(7) <= pprod(16) (19);
st7col53(7) <= pprod(16) (20);
st7col54(6) <= pprod(16) (21);
st7col55(6) <= pprod(16) (22);
st7col56(5) <= pprod(16) (23);
st7col57(5) <= pprod(16) (24);
st7col58(4) <= pprod(16) (25);
st7col59(4) <= pprod(16) (26);
st7col60(3) <= pprod(16) (27);
st7col61(3) <= pprod(16) (28);
st7col62(2) <= pprod(16) (29);
st7col63(2) <= pprod(16) (30);
st7col64(1) <= pprod(16) (31);
res_a <= st1col64(0) & st1col63(0) & st1col62(0) & st1col61(0) & st1col60(0) & st1col59(0) & st1col58(0) & st1col57(0) & st1col56(0) & st1col55(0) & st1col54(0) & st1col53(0) & st1col52(0) & st1col51(0) & st1col50(0) & st1col49(0) & st1col48(0) & st1col47(0) & st1col46(0) & st1col45(0) & st1col44(0) & st1col43(0) & st1col42(0) & st1col41(0) & st1col40(0) & st1col39(0) & st1col38(0) & st1col37(0) & st1col36(0) & st1col35(0) & st1col34(0) & st1col33(0) & st1col32(0) & st1col31(0) & st1col30(0) & st1col29(0) & st1col28(0) & st1col27(0) & st1col26(0) & st1col25(0) & st1col24(0) & st1col23(0) & st1col22(0) & st1col21(0) & st1col20(0) & st1col19(0) & st1col18(0) & st1col17(0) & st1col16(0) & st1col15(0) & st1col14(0) & st1col13(0) & st1col12(0) & st1col11(0) & st1col10(0) & st1col9(0) & st1col8(0) & st1col7(0) & st1col6(0) & st1col5(0) & st1col4(0) & st1col3(0) & st1col2(0) & st1col1(0);
res_b <= st1col64(1) & st1col63(1) & st1col62(1) & st1col61(1) & st1col60(1) & st1col59(1) & st1col58(1) & st1col57(1) & st1col56(1) & st1col55(1) & st1col54(1) & st1col53(1) & st1col52(1) & st1col51(1) & st1col50(1) & st1col49(1) & st1col48(1) & st1col47(1) & st1col46(1) & st1col45(1) & st1col44(1) & st1col43(1) & st1col42(1) & st1col41(1) & st1col40(1) & st1col39(1) & st1col38(1) & st1col37(1) & st1col36(1) & st1col35(1) & st1col34(1) & st1col33(1) & st1col32(1) & st1col31(1) & st1col30(1) & st1col29(1) & st1col28(1) & st1col27(1) & st1col26(1) & st1col25(1) & st1col24(1) & st1col23(1) & st1col22(1) & st1col21(1) & st1col20(1) & st1col19(1) & st1col18(1) & st1col17(1) & st1col16(1) & st1col15(1) & st1col14(1) & st1col13(1) & st1col12(1) & st1col11(1) & st1col10(1) & st1col9(1) & st1col8(1) & st1col7(1) & st1col6(1) & st1col5(1) & st1col4(1) & st1col3(1) & '0' & st1col1(1);

-- END AUTOGEN COMPS

z <= std_logic_vector(unsigned(res_a) + unsigned(res_b));
end RTL;