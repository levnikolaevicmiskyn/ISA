

package simconsts is
	constant NPIPE : integer := 1;
	constant FIXED_PIPE: integer := 5;
end simconsts;

package body simconsts is
end simconsts;
