

package simconsts is
	constant NPIPE : integer := 1;
	constant FIXED_PIPE: integer := 4;
end simconsts;

package body simconsts is
end simconsts;
