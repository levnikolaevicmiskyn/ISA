library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MBE is
	generic(N:integer := 4);
	port(
		m_and, m_ier: in std_logic_vector(N-1 downto 0);
		z: out std_logic_vector(2*N-1 downto 0)
		);
end entity MBE;

architecture RTL of MBE is

component FA is
port(a, b, cin: in std_logic;
	s, cout: out std_logic);
end component;

component HA is
port(a, b: in std_logic;
	s, cout: out std_logic);
end component;
type matype is array(N/2 downto 0) of std_logic_vector(N downto 0); -- N/2 operands
signal pprod: matype;
signal a, a2, a_neg, a2_neg: std_logic_vector(N downto 0);
signal S: std_logic_vector(N/2 downto 0);
signal res_a, res_b: std_logic_vector(2*N-1 downto 0); 
 
-- BEGIN AUTOGEN DECL
signal st1col1: std_logic_vector(2-1 downto 0);
signal st1col2: std_logic_vector(1-1 downto 0);
signal st1col3: std_logic_vector(2-1 downto 0);
signal st1col4: std_logic_vector(2-1 downto 0);
signal st1col5: std_logic_vector(2-1 downto 0);
signal st1col6: std_logic_vector(2-1 downto 0);
signal st1col7: std_logic_vector(2-1 downto 0);
signal st1col8: std_logic_vector(2-1 downto 0);
signal st1col9: std_logic_vector(2-1 downto 0);
signal st1col10: std_logic_vector(2-1 downto 0);
signal st1col11: std_logic_vector(2-1 downto 0);
signal st1col12: std_logic_vector(2-1 downto 0);
signal st1col13: std_logic_vector(2-1 downto 0);
signal st1col14: std_logic_vector(2-1 downto 0);
signal st1col15: std_logic_vector(2-1 downto 0);
signal st1col16: std_logic_vector(2-1 downto 0);
signal st1col17: std_logic_vector(2-1 downto 0);
signal st1col18: std_logic_vector(2-1 downto 0);
signal st1col19: std_logic_vector(2-1 downto 0);
signal st1col20: std_logic_vector(2-1 downto 0);
signal st1col21: std_logic_vector(2-1 downto 0);
signal st1col22: std_logic_vector(2-1 downto 0);
signal st1col23: std_logic_vector(2-1 downto 0);
signal st1col24: std_logic_vector(2-1 downto 0);
signal st1col25: std_logic_vector(2-1 downto 0);
signal st1col26: std_logic_vector(2-1 downto 0);
signal st1col27: std_logic_vector(2-1 downto 0);
signal st1col28: std_logic_vector(2-1 downto 0);
signal st1col29: std_logic_vector(2-1 downto 0);
signal st1col30: std_logic_vector(2-1 downto 0);
signal st1col31: std_logic_vector(2-1 downto 0);
signal st1col32: std_logic_vector(2-1 downto 0);
signal st1col33: std_logic_vector(2-1 downto 0);
signal st1col34: std_logic_vector(2-1 downto 0);
signal st1col35: std_logic_vector(2-1 downto 0);
signal st1col36: std_logic_vector(2-1 downto 0);
signal st1col37: std_logic_vector(2-1 downto 0);
signal st1col38: std_logic_vector(2-1 downto 0);
signal st1col39: std_logic_vector(2-1 downto 0);
signal st1col40: std_logic_vector(2-1 downto 0);
signal st1col41: std_logic_vector(2-1 downto 0);
signal st1col42: std_logic_vector(2-1 downto 0);
signal st1col43: std_logic_vector(2-1 downto 0);
signal st1col44: std_logic_vector(2-1 downto 0);
signal st1col45: std_logic_vector(2-1 downto 0);
signal st1col46: std_logic_vector(2-1 downto 0);
signal st1col47: std_logic_vector(2-1 downto 0);
signal st1col48: std_logic_vector(2-1 downto 0);
signal st2col1: std_logic_vector(2-1 downto 0);
signal st2col2: std_logic_vector(1-1 downto 0);
signal st2col3: std_logic_vector(3-1 downto 0);
signal st2col4: std_logic_vector(2-1 downto 0);
signal st2col5: std_logic_vector(3-1 downto 0);
signal st2col6: std_logic_vector(3-1 downto 0);
signal st2col7: std_logic_vector(3-1 downto 0);
signal st2col8: std_logic_vector(3-1 downto 0);
signal st2col9: std_logic_vector(3-1 downto 0);
signal st2col10: std_logic_vector(3-1 downto 0);
signal st2col11: std_logic_vector(3-1 downto 0);
signal st2col12: std_logic_vector(3-1 downto 0);
signal st2col13: std_logic_vector(3-1 downto 0);
signal st2col14: std_logic_vector(3-1 downto 0);
signal st2col15: std_logic_vector(3-1 downto 0);
signal st2col16: std_logic_vector(3-1 downto 0);
signal st2col17: std_logic_vector(3-1 downto 0);
signal st2col18: std_logic_vector(3-1 downto 0);
signal st2col19: std_logic_vector(3-1 downto 0);
signal st2col20: std_logic_vector(3-1 downto 0);
signal st2col21: std_logic_vector(3-1 downto 0);
signal st2col22: std_logic_vector(3-1 downto 0);
signal st2col23: std_logic_vector(3-1 downto 0);
signal st2col24: std_logic_vector(3-1 downto 0);
signal st2col25: std_logic_vector(3-1 downto 0);
signal st2col26: std_logic_vector(3-1 downto 0);
signal st2col27: std_logic_vector(3-1 downto 0);
signal st2col28: std_logic_vector(3-1 downto 0);
signal st2col29: std_logic_vector(3-1 downto 0);
signal st2col30: std_logic_vector(3-1 downto 0);
signal st2col31: std_logic_vector(3-1 downto 0);
signal st2col32: std_logic_vector(3-1 downto 0);
signal st2col33: std_logic_vector(3-1 downto 0);
signal st2col34: std_logic_vector(3-1 downto 0);
signal st2col35: std_logic_vector(3-1 downto 0);
signal st2col36: std_logic_vector(3-1 downto 0);
signal st2col37: std_logic_vector(3-1 downto 0);
signal st2col38: std_logic_vector(3-1 downto 0);
signal st2col39: std_logic_vector(3-1 downto 0);
signal st2col40: std_logic_vector(3-1 downto 0);
signal st2col41: std_logic_vector(3-1 downto 0);
signal st2col42: std_logic_vector(3-1 downto 0);
signal st2col43: std_logic_vector(3-1 downto 0);
signal st2col44: std_logic_vector(3-1 downto 0);
signal st2col45: std_logic_vector(3-1 downto 0);
signal st2col46: std_logic_vector(3-1 downto 0);
signal st2col47: std_logic_vector(3-1 downto 0);
signal st2col48: std_logic_vector(3-1 downto 0);
signal st3col1: std_logic_vector(2-1 downto 0);
signal st3col2: std_logic_vector(1-1 downto 0);
signal st3col3: std_logic_vector(3-1 downto 0);
signal st3col4: std_logic_vector(2-1 downto 0);
signal st3col5: std_logic_vector(4-1 downto 0);
signal st3col6: std_logic_vector(3-1 downto 0);
signal st3col7: std_logic_vector(4-1 downto 0);
signal st3col8: std_logic_vector(4-1 downto 0);
signal st3col9: std_logic_vector(4-1 downto 0);
signal st3col10: std_logic_vector(4-1 downto 0);
signal st3col11: std_logic_vector(4-1 downto 0);
signal st3col12: std_logic_vector(4-1 downto 0);
signal st3col13: std_logic_vector(4-1 downto 0);
signal st3col14: std_logic_vector(4-1 downto 0);
signal st3col15: std_logic_vector(4-1 downto 0);
signal st3col16: std_logic_vector(4-1 downto 0);
signal st3col17: std_logic_vector(4-1 downto 0);
signal st3col18: std_logic_vector(4-1 downto 0);
signal st3col19: std_logic_vector(4-1 downto 0);
signal st3col20: std_logic_vector(4-1 downto 0);
signal st3col21: std_logic_vector(4-1 downto 0);
signal st3col22: std_logic_vector(4-1 downto 0);
signal st3col23: std_logic_vector(4-1 downto 0);
signal st3col24: std_logic_vector(4-1 downto 0);
signal st3col25: std_logic_vector(4-1 downto 0);
signal st3col26: std_logic_vector(4-1 downto 0);
signal st3col27: std_logic_vector(4-1 downto 0);
signal st3col28: std_logic_vector(4-1 downto 0);
signal st3col29: std_logic_vector(4-1 downto 0);
signal st3col30: std_logic_vector(4-1 downto 0);
signal st3col31: std_logic_vector(4-1 downto 0);
signal st3col32: std_logic_vector(4-1 downto 0);
signal st3col33: std_logic_vector(4-1 downto 0);
signal st3col34: std_logic_vector(4-1 downto 0);
signal st3col35: std_logic_vector(4-1 downto 0);
signal st3col36: std_logic_vector(4-1 downto 0);
signal st3col37: std_logic_vector(4-1 downto 0);
signal st3col38: std_logic_vector(4-1 downto 0);
signal st3col39: std_logic_vector(4-1 downto 0);
signal st3col40: std_logic_vector(4-1 downto 0);
signal st3col41: std_logic_vector(4-1 downto 0);
signal st3col42: std_logic_vector(4-1 downto 0);
signal st3col43: std_logic_vector(4-1 downto 0);
signal st3col44: std_logic_vector(4-1 downto 0);
signal st3col45: std_logic_vector(4-1 downto 0);
signal st3col46: std_logic_vector(4-1 downto 0);
signal st3col47: std_logic_vector(3-1 downto 0);
signal st3col48: std_logic_vector(2-1 downto 0);
signal st4col1: std_logic_vector(2-1 downto 0);
signal st4col2: std_logic_vector(1-1 downto 0);
signal st4col3: std_logic_vector(3-1 downto 0);
signal st4col4: std_logic_vector(2-1 downto 0);
signal st4col5: std_logic_vector(4-1 downto 0);
signal st4col6: std_logic_vector(3-1 downto 0);
signal st4col7: std_logic_vector(5-1 downto 0);
signal st4col8: std_logic_vector(4-1 downto 0);
signal st4col9: std_logic_vector(6-1 downto 0);
signal st4col10: std_logic_vector(5-1 downto 0);
signal st4col11: std_logic_vector(6-1 downto 0);
signal st4col12: std_logic_vector(6-1 downto 0);
signal st4col13: std_logic_vector(6-1 downto 0);
signal st4col14: std_logic_vector(6-1 downto 0);
signal st4col15: std_logic_vector(6-1 downto 0);
signal st4col16: std_logic_vector(6-1 downto 0);
signal st4col17: std_logic_vector(6-1 downto 0);
signal st4col18: std_logic_vector(6-1 downto 0);
signal st4col19: std_logic_vector(6-1 downto 0);
signal st4col20: std_logic_vector(6-1 downto 0);
signal st4col21: std_logic_vector(6-1 downto 0);
signal st4col22: std_logic_vector(6-1 downto 0);
signal st4col23: std_logic_vector(6-1 downto 0);
signal st4col24: std_logic_vector(6-1 downto 0);
signal st4col25: std_logic_vector(6-1 downto 0);
signal st4col26: std_logic_vector(6-1 downto 0);
signal st4col27: std_logic_vector(6-1 downto 0);
signal st4col28: std_logic_vector(6-1 downto 0);
signal st4col29: std_logic_vector(6-1 downto 0);
signal st4col30: std_logic_vector(6-1 downto 0);
signal st4col31: std_logic_vector(6-1 downto 0);
signal st4col32: std_logic_vector(6-1 downto 0);
signal st4col33: std_logic_vector(6-1 downto 0);
signal st4col34: std_logic_vector(6-1 downto 0);
signal st4col35: std_logic_vector(6-1 downto 0);
signal st4col36: std_logic_vector(6-1 downto 0);
signal st4col37: std_logic_vector(6-1 downto 0);
signal st4col38: std_logic_vector(6-1 downto 0);
signal st4col39: std_logic_vector(6-1 downto 0);
signal st4col40: std_logic_vector(6-1 downto 0);
signal st4col41: std_logic_vector(6-1 downto 0);
signal st4col42: std_logic_vector(6-1 downto 0);
signal st4col43: std_logic_vector(5-1 downto 0);
signal st4col44: std_logic_vector(4-1 downto 0);
signal st4col45: std_logic_vector(4-1 downto 0);
signal st4col46: std_logic_vector(3-1 downto 0);
signal st4col47: std_logic_vector(3-1 downto 0);
signal st4col48: std_logic_vector(2-1 downto 0);
signal st5col1: std_logic_vector(2-1 downto 0);
signal st5col2: std_logic_vector(1-1 downto 0);
signal st5col3: std_logic_vector(3-1 downto 0);
signal st5col4: std_logic_vector(2-1 downto 0);
signal st5col5: std_logic_vector(4-1 downto 0);
signal st5col6: std_logic_vector(3-1 downto 0);
signal st5col7: std_logic_vector(5-1 downto 0);
signal st5col8: std_logic_vector(4-1 downto 0);
signal st5col9: std_logic_vector(6-1 downto 0);
signal st5col10: std_logic_vector(5-1 downto 0);
signal st5col11: std_logic_vector(7-1 downto 0);
signal st5col12: std_logic_vector(6-1 downto 0);
signal st5col13: std_logic_vector(8-1 downto 0);
signal st5col14: std_logic_vector(7-1 downto 0);
signal st5col15: std_logic_vector(9-1 downto 0);
signal st5col16: std_logic_vector(8-1 downto 0);
signal st5col17: std_logic_vector(9-1 downto 0);
signal st5col18: std_logic_vector(9-1 downto 0);
signal st5col19: std_logic_vector(9-1 downto 0);
signal st5col20: std_logic_vector(9-1 downto 0);
signal st5col21: std_logic_vector(9-1 downto 0);
signal st5col22: std_logic_vector(9-1 downto 0);
signal st5col23: std_logic_vector(9-1 downto 0);
signal st5col24: std_logic_vector(9-1 downto 0);
signal st5col25: std_logic_vector(9-1 downto 0);
signal st5col26: std_logic_vector(9-1 downto 0);
signal st5col27: std_logic_vector(9-1 downto 0);
signal st5col28: std_logic_vector(9-1 downto 0);
signal st5col29: std_logic_vector(9-1 downto 0);
signal st5col30: std_logic_vector(9-1 downto 0);
signal st5col31: std_logic_vector(9-1 downto 0);
signal st5col32: std_logic_vector(9-1 downto 0);
signal st5col33: std_logic_vector(9-1 downto 0);
signal st5col34: std_logic_vector(9-1 downto 0);
signal st5col35: std_logic_vector(9-1 downto 0);
signal st5col36: std_logic_vector(9-1 downto 0);
signal st5col37: std_logic_vector(8-1 downto 0);
signal st5col38: std_logic_vector(7-1 downto 0);
signal st5col39: std_logic_vector(7-1 downto 0);
signal st5col40: std_logic_vector(6-1 downto 0);
signal st5col41: std_logic_vector(6-1 downto 0);
signal st5col42: std_logic_vector(5-1 downto 0);
signal st5col43: std_logic_vector(5-1 downto 0);
signal st5col44: std_logic_vector(4-1 downto 0);
signal st5col45: std_logic_vector(4-1 downto 0);
signal st5col46: std_logic_vector(3-1 downto 0);
signal st5col47: std_logic_vector(3-1 downto 0);
signal st5col48: std_logic_vector(2-1 downto 0);
signal st6col1: std_logic_vector(2-1 downto 0);
signal st6col2: std_logic_vector(1-1 downto 0);
signal st6col3: std_logic_vector(3-1 downto 0);
signal st6col4: std_logic_vector(2-1 downto 0);
signal st6col5: std_logic_vector(4-1 downto 0);
signal st6col6: std_logic_vector(3-1 downto 0);
signal st6col7: std_logic_vector(5-1 downto 0);
signal st6col8: std_logic_vector(4-1 downto 0);
signal st6col9: std_logic_vector(6-1 downto 0);
signal st6col10: std_logic_vector(5-1 downto 0);
signal st6col11: std_logic_vector(7-1 downto 0);
signal st6col12: std_logic_vector(6-1 downto 0);
signal st6col13: std_logic_vector(8-1 downto 0);
signal st6col14: std_logic_vector(7-1 downto 0);
signal st6col15: std_logic_vector(9-1 downto 0);
signal st6col16: std_logic_vector(8-1 downto 0);
signal st6col17: std_logic_vector(10-1 downto 0);
signal st6col18: std_logic_vector(9-1 downto 0);
signal st6col19: std_logic_vector(11-1 downto 0);
signal st6col20: std_logic_vector(10-1 downto 0);
signal st6col21: std_logic_vector(12-1 downto 0);
signal st6col22: std_logic_vector(11-1 downto 0);
signal st6col23: std_logic_vector(13-1 downto 0);
signal st6col24: std_logic_vector(12-1 downto 0);
signal st6col25: std_logic_vector(13-1 downto 0);
signal st6col26: std_logic_vector(13-1 downto 0);
signal st6col27: std_logic_vector(13-1 downto 0);
signal st6col28: std_logic_vector(13-1 downto 0);
signal st6col29: std_logic_vector(12-1 downto 0);
signal st6col30: std_logic_vector(11-1 downto 0);
signal st6col31: std_logic_vector(11-1 downto 0);
signal st6col32: std_logic_vector(10-1 downto 0);
signal st6col33: std_logic_vector(10-1 downto 0);
signal st6col34: std_logic_vector(9-1 downto 0);
signal st6col35: std_logic_vector(9-1 downto 0);
signal st6col36: std_logic_vector(8-1 downto 0);
signal st6col37: std_logic_vector(8-1 downto 0);
signal st6col38: std_logic_vector(7-1 downto 0);
signal st6col39: std_logic_vector(7-1 downto 0);
signal st6col40: std_logic_vector(6-1 downto 0);
signal st6col41: std_logic_vector(6-1 downto 0);
signal st6col42: std_logic_vector(5-1 downto 0);
signal st6col43: std_logic_vector(5-1 downto 0);
signal st6col44: std_logic_vector(4-1 downto 0);
signal st6col45: std_logic_vector(4-1 downto 0);
signal st6col46: std_logic_vector(3-1 downto 0);
signal st6col47: std_logic_vector(3-1 downto 0);
signal st6col48: std_logic_vector(2-1 downto 0);
-- END AUTOGEN DECL

begin
-- Extend multiplicand
a <= '0' & m_and;
a_neg_proc: process (a)
			begin
				for i in a'range loop
					a_neg(i) <= not a(i);
				end loop;
			end process;
			
a2_neg_proc: process (a2)
			begin
				for i in a2'range loop
					a2_neg(i) <= not a2(i);
				end loop;
			end process;
			
-- a2 = multiplicand * 2
a2 <= m_and & '0';

benc_proc: process(a, a2, a_neg, a2_neg, m_and, m_ier)
variable window: std_logic_vector(2 downto 0);
begin
	for i in 0 to N/2 loop
		if i = 0 then
			window := m_ier(1 downto 0) & '0';
		elsif i = N/2 then
			window := "00" & m_ier(N-1);
		else
			window := m_ier(2*i+1 downto 2*i-1);
		end if;
		
		if window = "000" then
			pprod(i) <= (OTHERS => '0');
		elsif window = "001" or window = "010" then
			pprod(i) <= a;
		elsif window = "101" or window = "110" then
			pprod(i) <= a_neg;
		elsif window = "011" then
			pprod(i) <= a2;
		elsif window = "100" then
			pprod(i) <= a2_neg;
		else -- elseif window = "111" then
			pprod(i) <= (OTHERS => '1');
		end if;
		
	S(i) <= window(2);
	end loop;
end process;

-- BEGIN AUTOGEN COMPS
st5col1(0)<=st6col1(0);
st5col1(1)<=st6col1(1);
st5col2(0)<=st6col2(0);
st5col3(0)<=st6col3(0);
st5col3(1)<=st6col3(1);
st5col3(2)<=st6col3(2);
st5col4(0)<=st6col4(0);
st5col4(1)<=st6col4(1);
st5col5(0)<=st6col5(0);
st5col5(1)<=st6col5(1);
st5col5(2)<=st6col5(2);
st5col5(3)<=st6col5(3);
st5col6(0)<=st6col6(0);
st5col6(1)<=st6col6(1);
st5col6(2)<=st6col6(2);
st5col7(0)<=st6col7(0);
st5col7(1)<=st6col7(1);
st5col7(2)<=st6col7(2);
st5col7(3)<=st6col7(3);
st5col7(4)<=st6col7(4);
st5col8(0)<=st6col8(0);
st5col8(1)<=st6col8(1);
st5col8(2)<=st6col8(2);
st5col8(3)<=st6col8(3);
st5col9(0)<=st6col9(0);
st5col9(1)<=st6col9(1);
st5col9(2)<=st6col9(2);
st5col9(3)<=st6col9(3);
st5col9(4)<=st6col9(4);
st5col9(5)<=st6col9(5);
st5col10(0)<=st6col10(0);
st5col10(1)<=st6col10(1);
st5col10(2)<=st6col10(2);
st5col10(3)<=st6col10(3);
st5col10(4)<=st6col10(4);
st5col11(0)<=st6col11(0);
st5col11(1)<=st6col11(1);
st5col11(2)<=st6col11(2);
st5col11(3)<=st6col11(3);
st5col11(4)<=st6col11(4);
st5col11(5)<=st6col11(5);
st5col11(6)<=st6col11(6);
st5col12(0)<=st6col12(0);
st5col12(1)<=st6col12(1);
st5col12(2)<=st6col12(2);
st5col12(3)<=st6col12(3);
st5col12(4)<=st6col12(4);
st5col12(5)<=st6col12(5);
st5col13(0)<=st6col13(0);
st5col13(1)<=st6col13(1);
st5col13(2)<=st6col13(2);
st5col13(3)<=st6col13(3);
st5col13(4)<=st6col13(4);
st5col13(5)<=st6col13(5);
st5col13(6)<=st6col13(6);
st5col13(7)<=st6col13(7);
st5col14(0)<=st6col14(0);
st5col14(1)<=st6col14(1);
st5col14(2)<=st6col14(2);
st5col14(3)<=st6col14(3);
st5col14(4)<=st6col14(4);
st5col14(5)<=st6col14(5);
st5col14(6)<=st6col14(6);
st5col15(0)<=st6col15(0);
st5col15(1)<=st6col15(1);
st5col15(2)<=st6col15(2);
st5col15(3)<=st6col15(3);
st5col15(4)<=st6col15(4);
st5col15(5)<=st6col15(5);
st5col15(6)<=st6col15(6);
st5col15(7)<=st6col15(7);
st5col15(8)<=st6col15(8);
st5col16(0)<=st6col16(0);
st5col16(1)<=st6col16(1);
st5col16(2)<=st6col16(2);
st5col16(3)<=st6col16(3);
st5col16(4)<=st6col16(4);
st5col16(5)<=st6col16(5);
st5col16(6)<=st6col16(6);
st5col16(7)<=st6col16(7);
ha1st6col17: HA port map(st6col17(0),st6col17(1),st5col17(0),st5col18(0));
st5col17(1)<=st6col17(2);
st5col17(2)<=st6col17(3);
st5col17(3)<=st6col17(4);
st5col17(4)<=st6col17(5);
st5col17(5)<=st6col17(6);
st5col17(6)<=st6col17(7);
st5col17(7)<=st6col17(8);
st5col17(8)<=st6col17(9);
ha1st6col18: HA port map(st6col18(0),st6col18(1),st5col18(1),st5col19(0));
st5col18(2)<=st6col18(2);
st5col18(3)<=st6col18(3);
st5col18(4)<=st6col18(4);
st5col18(5)<=st6col18(5);
st5col18(6)<=st6col18(6);
st5col18(7)<=st6col18(7);
st5col18(8)<=st6col18(8);
fa0st6col19: FA port map(st6col19(0),st6col19(1),st6col19(2),st5col19(1),st5col20(0));
ha1st6col19: HA port map(st6col19(3),st6col19(4),st5col19(2),st5col20(1));
st5col19(3)<=st6col19(5);
st5col19(4)<=st6col19(6);
st5col19(5)<=st6col19(7);
st5col19(6)<=st6col19(8);
st5col19(7)<=st6col19(9);
st5col19(8)<=st6col19(10);
fa0st6col20: FA port map(st6col20(0),st6col20(1),st6col20(2),st5col20(2),st5col21(0));
ha1st6col20: HA port map(st6col20(3),st6col20(4),st5col20(3),st5col21(1));
st5col20(4)<=st6col20(5);
st5col20(5)<=st6col20(6);
st5col20(6)<=st6col20(7);
st5col20(7)<=st6col20(8);
st5col20(8)<=st6col20(9);
fa0st6col21: FA port map(st6col21(0),st6col21(1),st6col21(2),st5col21(2),st5col22(0));
fa1st6col21: FA port map(st6col21(3),st6col21(4),st6col21(5),st5col21(3),st5col22(1));
ha1st6col21: HA port map(st6col21(6),st6col21(7),st5col21(4),st5col22(2));
st5col21(5)<=st6col21(8);
st5col21(6)<=st6col21(9);
st5col21(7)<=st6col21(10);
st5col21(8)<=st6col21(11);
fa0st6col22: FA port map(st6col22(0),st6col22(1),st6col22(2),st5col22(3),st5col23(0));
fa1st6col22: FA port map(st6col22(3),st6col22(4),st6col22(5),st5col22(4),st5col23(1));
ha1st6col22: HA port map(st6col22(6),st6col22(7),st5col22(5),st5col23(2));
st5col22(6)<=st6col22(8);
st5col22(7)<=st6col22(9);
st5col22(8)<=st6col22(10);
fa0st6col23: FA port map(st6col23(0),st6col23(1),st6col23(2),st5col23(3),st5col24(0));
fa1st6col23: FA port map(st6col23(3),st6col23(4),st6col23(5),st5col23(4),st5col24(1));
fa2st6col23: FA port map(st6col23(6),st6col23(7),st6col23(8),st5col23(5),st5col24(2));
ha1st6col23: HA port map(st6col23(9),st6col23(10),st5col23(6),st5col24(3));
st5col23(7)<=st6col23(11);
st5col23(8)<=st6col23(12);
fa0st6col24: FA port map(st6col24(0),st6col24(1),st6col24(2),st5col24(4),st5col25(0));
fa1st6col24: FA port map(st6col24(3),st6col24(4),st6col24(5),st5col24(5),st5col25(1));
fa2st6col24: FA port map(st6col24(6),st6col24(7),st6col24(8),st5col24(6),st5col25(2));
ha1st6col24: HA port map(st6col24(9),st6col24(10),st5col24(7),st5col25(3));
st5col24(8)<=st6col24(11);
fa0st6col25: FA port map(st6col25(0),st6col25(1),st6col25(2),st5col25(4),st5col26(0));
fa1st6col25: FA port map(st6col25(3),st6col25(4),st6col25(5),st5col25(5),st5col26(1));
fa2st6col25: FA port map(st6col25(6),st6col25(7),st6col25(8),st5col25(6),st5col26(2));
fa3st6col25: FA port map(st6col25(9),st6col25(10),st6col25(11),st5col25(7),st5col26(3));
st5col25(8)<=st6col25(12);
fa0st6col26: FA port map(st6col26(0),st6col26(1),st6col26(2),st5col26(4),st5col27(0));
fa1st6col26: FA port map(st6col26(3),st6col26(4),st6col26(5),st5col26(5),st5col27(1));
fa2st6col26: FA port map(st6col26(6),st6col26(7),st6col26(8),st5col26(6),st5col27(2));
fa3st6col26: FA port map(st6col26(9),st6col26(10),st6col26(11),st5col26(7),st5col27(3));
st5col26(8)<=st6col26(12);
fa0st6col27: FA port map(st6col27(0),st6col27(1),st6col27(2),st5col27(4),st5col28(0));
fa1st6col27: FA port map(st6col27(3),st6col27(4),st6col27(5),st5col27(5),st5col28(1));
fa2st6col27: FA port map(st6col27(6),st6col27(7),st6col27(8),st5col27(6),st5col28(2));
fa3st6col27: FA port map(st6col27(9),st6col27(10),st6col27(11),st5col27(7),st5col28(3));
st5col27(8)<=st6col27(12);
fa0st6col28: FA port map(st6col28(0),st6col28(1),st6col28(2),st5col28(4),st5col29(0));
fa1st6col28: FA port map(st6col28(3),st6col28(4),st6col28(5),st5col28(5),st5col29(1));
fa2st6col28: FA port map(st6col28(6),st6col28(7),st6col28(8),st5col28(6),st5col29(2));
fa3st6col28: FA port map(st6col28(9),st6col28(10),st6col28(11),st5col28(7),st5col29(3));
st5col28(8)<=st6col28(12);
fa0st6col29: FA port map(st6col29(0),st6col29(1),st6col29(2),st5col29(4),st5col30(0));
fa1st6col29: FA port map(st6col29(3),st6col29(4),st6col29(5),st5col29(5),st5col30(1));
fa2st6col29: FA port map(st6col29(6),st6col29(7),st6col29(8),st5col29(6),st5col30(2));
ha1st6col29: HA port map(st6col29(9),st6col29(10),st5col29(7),st5col30(3));
st5col29(8)<=st6col29(11);
fa0st6col30: FA port map(st6col30(0),st6col30(1),st6col30(2),st5col30(4),st5col31(0));
fa1st6col30: FA port map(st6col30(3),st6col30(4),st6col30(5),st5col30(5),st5col31(1));
fa2st6col30: FA port map(st6col30(6),st6col30(7),st6col30(8),st5col30(6),st5col31(2));
st5col30(7)<=st6col30(9);
st5col30(8)<=st6col30(10);
fa0st6col31: FA port map(st6col31(0),st6col31(1),st6col31(2),st5col31(3),st5col32(0));
fa1st6col31: FA port map(st6col31(3),st6col31(4),st6col31(5),st5col31(4),st5col32(1));
ha1st6col31: HA port map(st6col31(6),st6col31(7),st5col31(5),st5col32(2));
st5col31(6)<=st6col31(8);
st5col31(7)<=st6col31(9);
st5col31(8)<=st6col31(10);
fa0st6col32: FA port map(st6col32(0),st6col32(1),st6col32(2),st5col32(3),st5col33(0));
fa1st6col32: FA port map(st6col32(3),st6col32(4),st6col32(5),st5col32(4),st5col33(1));
st5col32(5)<=st6col32(6);
st5col32(6)<=st6col32(7);
st5col32(7)<=st6col32(8);
st5col32(8)<=st6col32(9);
fa0st6col33: FA port map(st6col33(0),st6col33(1),st6col33(2),st5col33(2),st5col34(0));
ha1st6col33: HA port map(st6col33(3),st6col33(4),st5col33(3),st5col34(1));
st5col33(4)<=st6col33(5);
st5col33(5)<=st6col33(6);
st5col33(6)<=st6col33(7);
st5col33(7)<=st6col33(8);
st5col33(8)<=st6col33(9);
fa0st6col34: FA port map(st6col34(0),st6col34(1),st6col34(2),st5col34(2),st5col35(0));
st5col34(3)<=st6col34(3);
st5col34(4)<=st6col34(4);
st5col34(5)<=st6col34(5);
st5col34(6)<=st6col34(6);
st5col34(7)<=st6col34(7);
st5col34(8)<=st6col34(8);
ha1st6col35: HA port map(st6col35(0),st6col35(1),st5col35(1),st5col36(0));
st5col35(2)<=st6col35(2);
st5col35(3)<=st6col35(3);
st5col35(4)<=st6col35(4);
st5col35(5)<=st6col35(5);
st5col35(6)<=st6col35(6);
st5col35(7)<=st6col35(7);
st5col35(8)<=st6col35(8);
st5col36(1)<=st6col36(0);
st5col36(2)<=st6col36(1);
st5col36(3)<=st6col36(2);
st5col36(4)<=st6col36(3);
st5col36(5)<=st6col36(4);
st5col36(6)<=st6col36(5);
st5col36(7)<=st6col36(6);
st5col36(8)<=st6col36(7);
st5col37(0)<=st6col37(0);
st5col37(1)<=st6col37(1);
st5col37(2)<=st6col37(2);
st5col37(3)<=st6col37(3);
st5col37(4)<=st6col37(4);
st5col37(5)<=st6col37(5);
st5col37(6)<=st6col37(6);
st5col37(7)<=st6col37(7);
st5col38(0)<=st6col38(0);
st5col38(1)<=st6col38(1);
st5col38(2)<=st6col38(2);
st5col38(3)<=st6col38(3);
st5col38(4)<=st6col38(4);
st5col38(5)<=st6col38(5);
st5col38(6)<=st6col38(6);
st5col39(0)<=st6col39(0);
st5col39(1)<=st6col39(1);
st5col39(2)<=st6col39(2);
st5col39(3)<=st6col39(3);
st5col39(4)<=st6col39(4);
st5col39(5)<=st6col39(5);
st5col39(6)<=st6col39(6);
st5col40(0)<=st6col40(0);
st5col40(1)<=st6col40(1);
st5col40(2)<=st6col40(2);
st5col40(3)<=st6col40(3);
st5col40(4)<=st6col40(4);
st5col40(5)<=st6col40(5);
st5col41(0)<=st6col41(0);
st5col41(1)<=st6col41(1);
st5col41(2)<=st6col41(2);
st5col41(3)<=st6col41(3);
st5col41(4)<=st6col41(4);
st5col41(5)<=st6col41(5);
st5col42(0)<=st6col42(0);
st5col42(1)<=st6col42(1);
st5col42(2)<=st6col42(2);
st5col42(3)<=st6col42(3);
st5col42(4)<=st6col42(4);
st5col43(0)<=st6col43(0);
st5col43(1)<=st6col43(1);
st5col43(2)<=st6col43(2);
st5col43(3)<=st6col43(3);
st5col43(4)<=st6col43(4);
st5col44(0)<=st6col44(0);
st5col44(1)<=st6col44(1);
st5col44(2)<=st6col44(2);
st5col44(3)<=st6col44(3);
st5col45(0)<=st6col45(0);
st5col45(1)<=st6col45(1);
st5col45(2)<=st6col45(2);
st5col45(3)<=st6col45(3);
st5col46(0)<=st6col46(0);
st5col46(1)<=st6col46(1);
st5col46(2)<=st6col46(2);
st5col47(0)<=st6col47(0);
st5col47(1)<=st6col47(1);
st5col47(2)<=st6col47(2);
st5col48(0)<=st6col48(0);
st5col48(1)<=st6col48(1);
st4col1(0)<=st5col1(0);
st4col1(1)<=st5col1(1);
st4col2(0)<=st5col2(0);
st4col3(0)<=st5col3(0);
st4col3(1)<=st5col3(1);
st4col3(2)<=st5col3(2);
st4col4(0)<=st5col4(0);
st4col4(1)<=st5col4(1);
st4col5(0)<=st5col5(0);
st4col5(1)<=st5col5(1);
st4col5(2)<=st5col5(2);
st4col5(3)<=st5col5(3);
st4col6(0)<=st5col6(0);
st4col6(1)<=st5col6(1);
st4col6(2)<=st5col6(2);
st4col7(0)<=st5col7(0);
st4col7(1)<=st5col7(1);
st4col7(2)<=st5col7(2);
st4col7(3)<=st5col7(3);
st4col7(4)<=st5col7(4);
st4col8(0)<=st5col8(0);
st4col8(1)<=st5col8(1);
st4col8(2)<=st5col8(2);
st4col8(3)<=st5col8(3);
st4col9(0)<=st5col9(0);
st4col9(1)<=st5col9(1);
st4col9(2)<=st5col9(2);
st4col9(3)<=st5col9(3);
st4col9(4)<=st5col9(4);
st4col9(5)<=st5col9(5);
st4col10(0)<=st5col10(0);
st4col10(1)<=st5col10(1);
st4col10(2)<=st5col10(2);
st4col10(3)<=st5col10(3);
st4col10(4)<=st5col10(4);
ha1st5col11: HA port map(st5col11(0),st5col11(1),st4col11(0),st4col12(0));
st4col11(1)<=st5col11(2);
st4col11(2)<=st5col11(3);
st4col11(3)<=st5col11(4);
st4col11(4)<=st5col11(5);
st4col11(5)<=st5col11(6);
ha1st5col12: HA port map(st5col12(0),st5col12(1),st4col12(1),st4col13(0));
st4col12(2)<=st5col12(2);
st4col12(3)<=st5col12(3);
st4col12(4)<=st5col12(4);
st4col12(5)<=st5col12(5);
fa0st5col13: FA port map(st5col13(0),st5col13(1),st5col13(2),st4col13(1),st4col14(0));
ha1st5col13: HA port map(st5col13(3),st5col13(4),st4col13(2),st4col14(1));
st4col13(3)<=st5col13(5);
st4col13(4)<=st5col13(6);
st4col13(5)<=st5col13(7);
fa0st5col14: FA port map(st5col14(0),st5col14(1),st5col14(2),st4col14(2),st4col15(0));
ha1st5col14: HA port map(st5col14(3),st5col14(4),st4col14(3),st4col15(1));
st4col14(4)<=st5col14(5);
st4col14(5)<=st5col14(6);
fa0st5col15: FA port map(st5col15(0),st5col15(1),st5col15(2),st4col15(2),st4col16(0));
fa1st5col15: FA port map(st5col15(3),st5col15(4),st5col15(5),st4col15(3),st4col16(1));
ha1st5col15: HA port map(st5col15(6),st5col15(7),st4col15(4),st4col16(2));
st4col15(5)<=st5col15(8);
fa0st5col16: FA port map(st5col16(0),st5col16(1),st5col16(2),st4col16(3),st4col17(0));
fa1st5col16: FA port map(st5col16(3),st5col16(4),st5col16(5),st4col16(4),st4col17(1));
ha1st5col16: HA port map(st5col16(6),st5col16(7),st4col16(5),st4col17(2));
fa0st5col17: FA port map(st5col17(0),st5col17(1),st5col17(2),st4col17(3),st4col18(0));
fa1st5col17: FA port map(st5col17(3),st5col17(4),st5col17(5),st4col17(4),st4col18(1));
fa2st5col17: FA port map(st5col17(6),st5col17(7),st5col17(8),st4col17(5),st4col18(2));
fa0st5col18: FA port map(st5col18(0),st5col18(1),st5col18(2),st4col18(3),st4col19(0));
fa1st5col18: FA port map(st5col18(3),st5col18(4),st5col18(5),st4col18(4),st4col19(1));
fa2st5col18: FA port map(st5col18(6),st5col18(7),st5col18(8),st4col18(5),st4col19(2));
fa0st5col19: FA port map(st5col19(0),st5col19(1),st5col19(2),st4col19(3),st4col20(0));
fa1st5col19: FA port map(st5col19(3),st5col19(4),st5col19(5),st4col19(4),st4col20(1));
fa2st5col19: FA port map(st5col19(6),st5col19(7),st5col19(8),st4col19(5),st4col20(2));
fa0st5col20: FA port map(st5col20(0),st5col20(1),st5col20(2),st4col20(3),st4col21(0));
fa1st5col20: FA port map(st5col20(3),st5col20(4),st5col20(5),st4col20(4),st4col21(1));
fa2st5col20: FA port map(st5col20(6),st5col20(7),st5col20(8),st4col20(5),st4col21(2));
fa0st5col21: FA port map(st5col21(0),st5col21(1),st5col21(2),st4col21(3),st4col22(0));
fa1st5col21: FA port map(st5col21(3),st5col21(4),st5col21(5),st4col21(4),st4col22(1));
fa2st5col21: FA port map(st5col21(6),st5col21(7),st5col21(8),st4col21(5),st4col22(2));
fa0st5col22: FA port map(st5col22(0),st5col22(1),st5col22(2),st4col22(3),st4col23(0));
fa1st5col22: FA port map(st5col22(3),st5col22(4),st5col22(5),st4col22(4),st4col23(1));
fa2st5col22: FA port map(st5col22(6),st5col22(7),st5col22(8),st4col22(5),st4col23(2));
fa0st5col23: FA port map(st5col23(0),st5col23(1),st5col23(2),st4col23(3),st4col24(0));
fa1st5col23: FA port map(st5col23(3),st5col23(4),st5col23(5),st4col23(4),st4col24(1));
fa2st5col23: FA port map(st5col23(6),st5col23(7),st5col23(8),st4col23(5),st4col24(2));
fa0st5col24: FA port map(st5col24(0),st5col24(1),st5col24(2),st4col24(3),st4col25(0));
fa1st5col24: FA port map(st5col24(3),st5col24(4),st5col24(5),st4col24(4),st4col25(1));
fa2st5col24: FA port map(st5col24(6),st5col24(7),st5col24(8),st4col24(5),st4col25(2));
fa0st5col25: FA port map(st5col25(0),st5col25(1),st5col25(2),st4col25(3),st4col26(0));
fa1st5col25: FA port map(st5col25(3),st5col25(4),st5col25(5),st4col25(4),st4col26(1));
fa2st5col25: FA port map(st5col25(6),st5col25(7),st5col25(8),st4col25(5),st4col26(2));
fa0st5col26: FA port map(st5col26(0),st5col26(1),st5col26(2),st4col26(3),st4col27(0));
fa1st5col26: FA port map(st5col26(3),st5col26(4),st5col26(5),st4col26(4),st4col27(1));
fa2st5col26: FA port map(st5col26(6),st5col26(7),st5col26(8),st4col26(5),st4col27(2));
fa0st5col27: FA port map(st5col27(0),st5col27(1),st5col27(2),st4col27(3),st4col28(0));
fa1st5col27: FA port map(st5col27(3),st5col27(4),st5col27(5),st4col27(4),st4col28(1));
fa2st5col27: FA port map(st5col27(6),st5col27(7),st5col27(8),st4col27(5),st4col28(2));
fa0st5col28: FA port map(st5col28(0),st5col28(1),st5col28(2),st4col28(3),st4col29(0));
fa1st5col28: FA port map(st5col28(3),st5col28(4),st5col28(5),st4col28(4),st4col29(1));
fa2st5col28: FA port map(st5col28(6),st5col28(7),st5col28(8),st4col28(5),st4col29(2));
fa0st5col29: FA port map(st5col29(0),st5col29(1),st5col29(2),st4col29(3),st4col30(0));
fa1st5col29: FA port map(st5col29(3),st5col29(4),st5col29(5),st4col29(4),st4col30(1));
fa2st5col29: FA port map(st5col29(6),st5col29(7),st5col29(8),st4col29(5),st4col30(2));
fa0st5col30: FA port map(st5col30(0),st5col30(1),st5col30(2),st4col30(3),st4col31(0));
fa1st5col30: FA port map(st5col30(3),st5col30(4),st5col30(5),st4col30(4),st4col31(1));
fa2st5col30: FA port map(st5col30(6),st5col30(7),st5col30(8),st4col30(5),st4col31(2));
fa0st5col31: FA port map(st5col31(0),st5col31(1),st5col31(2),st4col31(3),st4col32(0));
fa1st5col31: FA port map(st5col31(3),st5col31(4),st5col31(5),st4col31(4),st4col32(1));
fa2st5col31: FA port map(st5col31(6),st5col31(7),st5col31(8),st4col31(5),st4col32(2));
fa0st5col32: FA port map(st5col32(0),st5col32(1),st5col32(2),st4col32(3),st4col33(0));
fa1st5col32: FA port map(st5col32(3),st5col32(4),st5col32(5),st4col32(4),st4col33(1));
fa2st5col32: FA port map(st5col32(6),st5col32(7),st5col32(8),st4col32(5),st4col33(2));
fa0st5col33: FA port map(st5col33(0),st5col33(1),st5col33(2),st4col33(3),st4col34(0));
fa1st5col33: FA port map(st5col33(3),st5col33(4),st5col33(5),st4col33(4),st4col34(1));
fa2st5col33: FA port map(st5col33(6),st5col33(7),st5col33(8),st4col33(5),st4col34(2));
fa0st5col34: FA port map(st5col34(0),st5col34(1),st5col34(2),st4col34(3),st4col35(0));
fa1st5col34: FA port map(st5col34(3),st5col34(4),st5col34(5),st4col34(4),st4col35(1));
fa2st5col34: FA port map(st5col34(6),st5col34(7),st5col34(8),st4col34(5),st4col35(2));
fa0st5col35: FA port map(st5col35(0),st5col35(1),st5col35(2),st4col35(3),st4col36(0));
fa1st5col35: FA port map(st5col35(3),st5col35(4),st5col35(5),st4col35(4),st4col36(1));
fa2st5col35: FA port map(st5col35(6),st5col35(7),st5col35(8),st4col35(5),st4col36(2));
fa0st5col36: FA port map(st5col36(0),st5col36(1),st5col36(2),st4col36(3),st4col37(0));
fa1st5col36: FA port map(st5col36(3),st5col36(4),st5col36(5),st4col36(4),st4col37(1));
fa2st5col36: FA port map(st5col36(6),st5col36(7),st5col36(8),st4col36(5),st4col37(2));
fa0st5col37: FA port map(st5col37(0),st5col37(1),st5col37(2),st4col37(3),st4col38(0));
fa1st5col37: FA port map(st5col37(3),st5col37(4),st5col37(5),st4col37(4),st4col38(1));
ha1st5col37: HA port map(st5col37(6),st5col37(7),st4col37(5),st4col38(2));
fa0st5col38: FA port map(st5col38(0),st5col38(1),st5col38(2),st4col38(3),st4col39(0));
fa1st5col38: FA port map(st5col38(3),st5col38(4),st5col38(5),st4col38(4),st4col39(1));
st4col38(5)<=st5col38(6);
fa0st5col39: FA port map(st5col39(0),st5col39(1),st5col39(2),st4col39(2),st4col40(0));
ha1st5col39: HA port map(st5col39(3),st5col39(4),st4col39(3),st4col40(1));
st4col39(4)<=st5col39(5);
st4col39(5)<=st5col39(6);
fa0st5col40: FA port map(st5col40(0),st5col40(1),st5col40(2),st4col40(2),st4col41(0));
st4col40(3)<=st5col40(3);
st4col40(4)<=st5col40(4);
st4col40(5)<=st5col40(5);
ha1st5col41: HA port map(st5col41(0),st5col41(1),st4col41(1),st4col42(0));
st4col41(2)<=st5col41(2);
st4col41(3)<=st5col41(3);
st4col41(4)<=st5col41(4);
st4col41(5)<=st5col41(5);
st4col42(1)<=st5col42(0);
st4col42(2)<=st5col42(1);
st4col42(3)<=st5col42(2);
st4col42(4)<=st5col42(3);
st4col42(5)<=st5col42(4);
st4col43(0)<=st5col43(0);
st4col43(1)<=st5col43(1);
st4col43(2)<=st5col43(2);
st4col43(3)<=st5col43(3);
st4col43(4)<=st5col43(4);
st4col44(0)<=st5col44(0);
st4col44(1)<=st5col44(1);
st4col44(2)<=st5col44(2);
st4col44(3)<=st5col44(3);
st4col45(0)<=st5col45(0);
st4col45(1)<=st5col45(1);
st4col45(2)<=st5col45(2);
st4col45(3)<=st5col45(3);
st4col46(0)<=st5col46(0);
st4col46(1)<=st5col46(1);
st4col46(2)<=st5col46(2);
st4col47(0)<=st5col47(0);
st4col47(1)<=st5col47(1);
st4col47(2)<=st5col47(2);
st4col48(0)<=st5col48(0);
st4col48(1)<=st5col48(1);
st3col1(0)<=st4col1(0);
st3col1(1)<=st4col1(1);
st3col2(0)<=st4col2(0);
st3col3(0)<=st4col3(0);
st3col3(1)<=st4col3(1);
st3col3(2)<=st4col3(2);
st3col4(0)<=st4col4(0);
st3col4(1)<=st4col4(1);
st3col5(0)<=st4col5(0);
st3col5(1)<=st4col5(1);
st3col5(2)<=st4col5(2);
st3col5(3)<=st4col5(3);
st3col6(0)<=st4col6(0);
st3col6(1)<=st4col6(1);
st3col6(2)<=st4col6(2);
ha1st4col7: HA port map(st4col7(0),st4col7(1),st3col7(0),st3col8(0));
st3col7(1)<=st4col7(2);
st3col7(2)<=st4col7(3);
st3col7(3)<=st4col7(4);
ha1st4col8: HA port map(st4col8(0),st4col8(1),st3col8(1),st3col9(0));
st3col8(2)<=st4col8(2);
st3col8(3)<=st4col8(3);
fa0st4col9: FA port map(st4col9(0),st4col9(1),st4col9(2),st3col9(1),st3col10(0));
ha1st4col9: HA port map(st4col9(3),st4col9(4),st3col9(2),st3col10(1));
st3col9(3)<=st4col9(5);
fa0st4col10: FA port map(st4col10(0),st4col10(1),st4col10(2),st3col10(2),st3col11(0));
ha1st4col10: HA port map(st4col10(3),st4col10(4),st3col10(3),st3col11(1));
fa0st4col11: FA port map(st4col11(0),st4col11(1),st4col11(2),st3col11(2),st3col12(0));
fa1st4col11: FA port map(st4col11(3),st4col11(4),st4col11(5),st3col11(3),st3col12(1));
fa0st4col12: FA port map(st4col12(0),st4col12(1),st4col12(2),st3col12(2),st3col13(0));
fa1st4col12: FA port map(st4col12(3),st4col12(4),st4col12(5),st3col12(3),st3col13(1));
fa0st4col13: FA port map(st4col13(0),st4col13(1),st4col13(2),st3col13(2),st3col14(0));
fa1st4col13: FA port map(st4col13(3),st4col13(4),st4col13(5),st3col13(3),st3col14(1));
fa0st4col14: FA port map(st4col14(0),st4col14(1),st4col14(2),st3col14(2),st3col15(0));
fa1st4col14: FA port map(st4col14(3),st4col14(4),st4col14(5),st3col14(3),st3col15(1));
fa0st4col15: FA port map(st4col15(0),st4col15(1),st4col15(2),st3col15(2),st3col16(0));
fa1st4col15: FA port map(st4col15(3),st4col15(4),st4col15(5),st3col15(3),st3col16(1));
fa0st4col16: FA port map(st4col16(0),st4col16(1),st4col16(2),st3col16(2),st3col17(0));
fa1st4col16: FA port map(st4col16(3),st4col16(4),st4col16(5),st3col16(3),st3col17(1));
fa0st4col17: FA port map(st4col17(0),st4col17(1),st4col17(2),st3col17(2),st3col18(0));
fa1st4col17: FA port map(st4col17(3),st4col17(4),st4col17(5),st3col17(3),st3col18(1));
fa0st4col18: FA port map(st4col18(0),st4col18(1),st4col18(2),st3col18(2),st3col19(0));
fa1st4col18: FA port map(st4col18(3),st4col18(4),st4col18(5),st3col18(3),st3col19(1));
fa0st4col19: FA port map(st4col19(0),st4col19(1),st4col19(2),st3col19(2),st3col20(0));
fa1st4col19: FA port map(st4col19(3),st4col19(4),st4col19(5),st3col19(3),st3col20(1));
fa0st4col20: FA port map(st4col20(0),st4col20(1),st4col20(2),st3col20(2),st3col21(0));
fa1st4col20: FA port map(st4col20(3),st4col20(4),st4col20(5),st3col20(3),st3col21(1));
fa0st4col21: FA port map(st4col21(0),st4col21(1),st4col21(2),st3col21(2),st3col22(0));
fa1st4col21: FA port map(st4col21(3),st4col21(4),st4col21(5),st3col21(3),st3col22(1));
fa0st4col22: FA port map(st4col22(0),st4col22(1),st4col22(2),st3col22(2),st3col23(0));
fa1st4col22: FA port map(st4col22(3),st4col22(4),st4col22(5),st3col22(3),st3col23(1));
fa0st4col23: FA port map(st4col23(0),st4col23(1),st4col23(2),st3col23(2),st3col24(0));
fa1st4col23: FA port map(st4col23(3),st4col23(4),st4col23(5),st3col23(3),st3col24(1));
fa0st4col24: FA port map(st4col24(0),st4col24(1),st4col24(2),st3col24(2),st3col25(0));
fa1st4col24: FA port map(st4col24(3),st4col24(4),st4col24(5),st3col24(3),st3col25(1));
fa0st4col25: FA port map(st4col25(0),st4col25(1),st4col25(2),st3col25(2),st3col26(0));
fa1st4col25: FA port map(st4col25(3),st4col25(4),st4col25(5),st3col25(3),st3col26(1));
fa0st4col26: FA port map(st4col26(0),st4col26(1),st4col26(2),st3col26(2),st3col27(0));
fa1st4col26: FA port map(st4col26(3),st4col26(4),st4col26(5),st3col26(3),st3col27(1));
fa0st4col27: FA port map(st4col27(0),st4col27(1),st4col27(2),st3col27(2),st3col28(0));
fa1st4col27: FA port map(st4col27(3),st4col27(4),st4col27(5),st3col27(3),st3col28(1));
fa0st4col28: FA port map(st4col28(0),st4col28(1),st4col28(2),st3col28(2),st3col29(0));
fa1st4col28: FA port map(st4col28(3),st4col28(4),st4col28(5),st3col28(3),st3col29(1));
fa0st4col29: FA port map(st4col29(0),st4col29(1),st4col29(2),st3col29(2),st3col30(0));
fa1st4col29: FA port map(st4col29(3),st4col29(4),st4col29(5),st3col29(3),st3col30(1));
fa0st4col30: FA port map(st4col30(0),st4col30(1),st4col30(2),st3col30(2),st3col31(0));
fa1st4col30: FA port map(st4col30(3),st4col30(4),st4col30(5),st3col30(3),st3col31(1));
fa0st4col31: FA port map(st4col31(0),st4col31(1),st4col31(2),st3col31(2),st3col32(0));
fa1st4col31: FA port map(st4col31(3),st4col31(4),st4col31(5),st3col31(3),st3col32(1));
fa0st4col32: FA port map(st4col32(0),st4col32(1),st4col32(2),st3col32(2),st3col33(0));
fa1st4col32: FA port map(st4col32(3),st4col32(4),st4col32(5),st3col32(3),st3col33(1));
fa0st4col33: FA port map(st4col33(0),st4col33(1),st4col33(2),st3col33(2),st3col34(0));
fa1st4col33: FA port map(st4col33(3),st4col33(4),st4col33(5),st3col33(3),st3col34(1));
fa0st4col34: FA port map(st4col34(0),st4col34(1),st4col34(2),st3col34(2),st3col35(0));
fa1st4col34: FA port map(st4col34(3),st4col34(4),st4col34(5),st3col34(3),st3col35(1));
fa0st4col35: FA port map(st4col35(0),st4col35(1),st4col35(2),st3col35(2),st3col36(0));
fa1st4col35: FA port map(st4col35(3),st4col35(4),st4col35(5),st3col35(3),st3col36(1));
fa0st4col36: FA port map(st4col36(0),st4col36(1),st4col36(2),st3col36(2),st3col37(0));
fa1st4col36: FA port map(st4col36(3),st4col36(4),st4col36(5),st3col36(3),st3col37(1));
fa0st4col37: FA port map(st4col37(0),st4col37(1),st4col37(2),st3col37(2),st3col38(0));
fa1st4col37: FA port map(st4col37(3),st4col37(4),st4col37(5),st3col37(3),st3col38(1));
fa0st4col38: FA port map(st4col38(0),st4col38(1),st4col38(2),st3col38(2),st3col39(0));
fa1st4col38: FA port map(st4col38(3),st4col38(4),st4col38(5),st3col38(3),st3col39(1));
fa0st4col39: FA port map(st4col39(0),st4col39(1),st4col39(2),st3col39(2),st3col40(0));
fa1st4col39: FA port map(st4col39(3),st4col39(4),st4col39(5),st3col39(3),st3col40(1));
fa0st4col40: FA port map(st4col40(0),st4col40(1),st4col40(2),st3col40(2),st3col41(0));
fa1st4col40: FA port map(st4col40(3),st4col40(4),st4col40(5),st3col40(3),st3col41(1));
fa0st4col41: FA port map(st4col41(0),st4col41(1),st4col41(2),st3col41(2),st3col42(0));
fa1st4col41: FA port map(st4col41(3),st4col41(4),st4col41(5),st3col41(3),st3col42(1));
fa0st4col42: FA port map(st4col42(0),st4col42(1),st4col42(2),st3col42(2),st3col43(0));
fa1st4col42: FA port map(st4col42(3),st4col42(4),st4col42(5),st3col42(3),st3col43(1));
fa0st4col43: FA port map(st4col43(0),st4col43(1),st4col43(2),st3col43(2),st3col44(0));
ha1st4col43: HA port map(st4col43(3),st4col43(4),st3col43(3),st3col44(1));
fa0st4col44: FA port map(st4col44(0),st4col44(1),st4col44(2),st3col44(2),st3col45(0));
st3col44(3)<=st4col44(3);
ha1st4col45: HA port map(st4col45(0),st4col45(1),st3col45(1),st3col46(0));
st3col45(2)<=st4col45(2);
st3col45(3)<=st4col45(3);
st3col46(1)<=st4col46(0);
st3col46(2)<=st4col46(1);
st3col46(3)<=st4col46(2);
st3col47(0)<=st4col47(0);
st3col47(1)<=st4col47(1);
st3col47(2)<=st4col47(2);
st3col48(0)<=st4col48(0);
st3col48(1)<=st4col48(1);
st2col1(0)<=st3col1(0);
st2col1(1)<=st3col1(1);
st2col2(0)<=st3col2(0);
st2col3(0)<=st3col3(0);
st2col3(1)<=st3col3(1);
st2col3(2)<=st3col3(2);
st2col4(0)<=st3col4(0);
st2col4(1)<=st3col4(1);
ha1st3col5: HA port map(st3col5(0),st3col5(1),st2col5(0),st2col6(0));
st2col5(1)<=st3col5(2);
st2col5(2)<=st3col5(3);
ha1st3col6: HA port map(st3col6(0),st3col6(1),st2col6(1),st2col7(0));
st2col6(2)<=st3col6(2);
fa0st3col7: FA port map(st3col7(0),st3col7(1),st3col7(2),st2col7(1),st2col8(0));
st2col7(2)<=st3col7(3);
fa0st3col8: FA port map(st3col8(0),st3col8(1),st3col8(2),st2col8(1),st2col9(0));
st2col8(2)<=st3col8(3);
fa0st3col9: FA port map(st3col9(0),st3col9(1),st3col9(2),st2col9(1),st2col10(0));
st2col9(2)<=st3col9(3);
fa0st3col10: FA port map(st3col10(0),st3col10(1),st3col10(2),st2col10(1),st2col11(0));
st2col10(2)<=st3col10(3);
fa0st3col11: FA port map(st3col11(0),st3col11(1),st3col11(2),st2col11(1),st2col12(0));
st2col11(2)<=st3col11(3);
fa0st3col12: FA port map(st3col12(0),st3col12(1),st3col12(2),st2col12(1),st2col13(0));
st2col12(2)<=st3col12(3);
fa0st3col13: FA port map(st3col13(0),st3col13(1),st3col13(2),st2col13(1),st2col14(0));
st2col13(2)<=st3col13(3);
fa0st3col14: FA port map(st3col14(0),st3col14(1),st3col14(2),st2col14(1),st2col15(0));
st2col14(2)<=st3col14(3);
fa0st3col15: FA port map(st3col15(0),st3col15(1),st3col15(2),st2col15(1),st2col16(0));
st2col15(2)<=st3col15(3);
fa0st3col16: FA port map(st3col16(0),st3col16(1),st3col16(2),st2col16(1),st2col17(0));
st2col16(2)<=st3col16(3);
fa0st3col17: FA port map(st3col17(0),st3col17(1),st3col17(2),st2col17(1),st2col18(0));
st2col17(2)<=st3col17(3);
fa0st3col18: FA port map(st3col18(0),st3col18(1),st3col18(2),st2col18(1),st2col19(0));
st2col18(2)<=st3col18(3);
fa0st3col19: FA port map(st3col19(0),st3col19(1),st3col19(2),st2col19(1),st2col20(0));
st2col19(2)<=st3col19(3);
fa0st3col20: FA port map(st3col20(0),st3col20(1),st3col20(2),st2col20(1),st2col21(0));
st2col20(2)<=st3col20(3);
fa0st3col21: FA port map(st3col21(0),st3col21(1),st3col21(2),st2col21(1),st2col22(0));
st2col21(2)<=st3col21(3);
fa0st3col22: FA port map(st3col22(0),st3col22(1),st3col22(2),st2col22(1),st2col23(0));
st2col22(2)<=st3col22(3);
fa0st3col23: FA port map(st3col23(0),st3col23(1),st3col23(2),st2col23(1),st2col24(0));
st2col23(2)<=st3col23(3);
fa0st3col24: FA port map(st3col24(0),st3col24(1),st3col24(2),st2col24(1),st2col25(0));
st2col24(2)<=st3col24(3);
fa0st3col25: FA port map(st3col25(0),st3col25(1),st3col25(2),st2col25(1),st2col26(0));
st2col25(2)<=st3col25(3);
fa0st3col26: FA port map(st3col26(0),st3col26(1),st3col26(2),st2col26(1),st2col27(0));
st2col26(2)<=st3col26(3);
fa0st3col27: FA port map(st3col27(0),st3col27(1),st3col27(2),st2col27(1),st2col28(0));
st2col27(2)<=st3col27(3);
fa0st3col28: FA port map(st3col28(0),st3col28(1),st3col28(2),st2col28(1),st2col29(0));
st2col28(2)<=st3col28(3);
fa0st3col29: FA port map(st3col29(0),st3col29(1),st3col29(2),st2col29(1),st2col30(0));
st2col29(2)<=st3col29(3);
fa0st3col30: FA port map(st3col30(0),st3col30(1),st3col30(2),st2col30(1),st2col31(0));
st2col30(2)<=st3col30(3);
fa0st3col31: FA port map(st3col31(0),st3col31(1),st3col31(2),st2col31(1),st2col32(0));
st2col31(2)<=st3col31(3);
fa0st3col32: FA port map(st3col32(0),st3col32(1),st3col32(2),st2col32(1),st2col33(0));
st2col32(2)<=st3col32(3);
fa0st3col33: FA port map(st3col33(0),st3col33(1),st3col33(2),st2col33(1),st2col34(0));
st2col33(2)<=st3col33(3);
fa0st3col34: FA port map(st3col34(0),st3col34(1),st3col34(2),st2col34(1),st2col35(0));
st2col34(2)<=st3col34(3);
fa0st3col35: FA port map(st3col35(0),st3col35(1),st3col35(2),st2col35(1),st2col36(0));
st2col35(2)<=st3col35(3);
fa0st3col36: FA port map(st3col36(0),st3col36(1),st3col36(2),st2col36(1),st2col37(0));
st2col36(2)<=st3col36(3);
fa0st3col37: FA port map(st3col37(0),st3col37(1),st3col37(2),st2col37(1),st2col38(0));
st2col37(2)<=st3col37(3);
fa0st3col38: FA port map(st3col38(0),st3col38(1),st3col38(2),st2col38(1),st2col39(0));
st2col38(2)<=st3col38(3);
fa0st3col39: FA port map(st3col39(0),st3col39(1),st3col39(2),st2col39(1),st2col40(0));
st2col39(2)<=st3col39(3);
fa0st3col40: FA port map(st3col40(0),st3col40(1),st3col40(2),st2col40(1),st2col41(0));
st2col40(2)<=st3col40(3);
fa0st3col41: FA port map(st3col41(0),st3col41(1),st3col41(2),st2col41(1),st2col42(0));
st2col41(2)<=st3col41(3);
fa0st3col42: FA port map(st3col42(0),st3col42(1),st3col42(2),st2col42(1),st2col43(0));
st2col42(2)<=st3col42(3);
fa0st3col43: FA port map(st3col43(0),st3col43(1),st3col43(2),st2col43(1),st2col44(0));
st2col43(2)<=st3col43(3);
fa0st3col44: FA port map(st3col44(0),st3col44(1),st3col44(2),st2col44(1),st2col45(0));
st2col44(2)<=st3col44(3);
fa0st3col45: FA port map(st3col45(0),st3col45(1),st3col45(2),st2col45(1),st2col46(0));
st2col45(2)<=st3col45(3);
fa0st3col46: FA port map(st3col46(0),st3col46(1),st3col46(2),st2col46(1),st2col47(0));
st2col46(2)<=st3col46(3);
ha1st3col47: HA port map(st3col47(0),st3col47(1),st2col47(1),st2col48(0));
st2col47(2)<=st3col47(2);
st2col48(1)<=st3col48(0);
st2col48(2)<=st3col48(1);
st1col1(0)<=st2col1(0);
st1col1(1)<=st2col1(1);
st1col2(0)<=st2col2(0);
ha1st2col3: HA port map(st2col3(0),st2col3(1),st1col3(0),st1col4(0));
st1col3(1)<=st2col3(2);
ha1st2col4: HA port map(st2col4(0),st2col4(1),st1col4(1),st1col5(0));
fa0st2col5: FA port map(st2col5(0),st2col5(1),st2col5(2),st1col5(1),st1col6(0));
fa0st2col6: FA port map(st2col6(0),st2col6(1),st2col6(2),st1col6(1),st1col7(0));
fa0st2col7: FA port map(st2col7(0),st2col7(1),st2col7(2),st1col7(1),st1col8(0));
fa0st2col8: FA port map(st2col8(0),st2col8(1),st2col8(2),st1col8(1),st1col9(0));
fa0st2col9: FA port map(st2col9(0),st2col9(1),st2col9(2),st1col9(1),st1col10(0));
fa0st2col10: FA port map(st2col10(0),st2col10(1),st2col10(2),st1col10(1),st1col11(0));
fa0st2col11: FA port map(st2col11(0),st2col11(1),st2col11(2),st1col11(1),st1col12(0));
fa0st2col12: FA port map(st2col12(0),st2col12(1),st2col12(2),st1col12(1),st1col13(0));
fa0st2col13: FA port map(st2col13(0),st2col13(1),st2col13(2),st1col13(1),st1col14(0));
fa0st2col14: FA port map(st2col14(0),st2col14(1),st2col14(2),st1col14(1),st1col15(0));
fa0st2col15: FA port map(st2col15(0),st2col15(1),st2col15(2),st1col15(1),st1col16(0));
fa0st2col16: FA port map(st2col16(0),st2col16(1),st2col16(2),st1col16(1),st1col17(0));
fa0st2col17: FA port map(st2col17(0),st2col17(1),st2col17(2),st1col17(1),st1col18(0));
fa0st2col18: FA port map(st2col18(0),st2col18(1),st2col18(2),st1col18(1),st1col19(0));
fa0st2col19: FA port map(st2col19(0),st2col19(1),st2col19(2),st1col19(1),st1col20(0));
fa0st2col20: FA port map(st2col20(0),st2col20(1),st2col20(2),st1col20(1),st1col21(0));
fa0st2col21: FA port map(st2col21(0),st2col21(1),st2col21(2),st1col21(1),st1col22(0));
fa0st2col22: FA port map(st2col22(0),st2col22(1),st2col22(2),st1col22(1),st1col23(0));
fa0st2col23: FA port map(st2col23(0),st2col23(1),st2col23(2),st1col23(1),st1col24(0));
fa0st2col24: FA port map(st2col24(0),st2col24(1),st2col24(2),st1col24(1),st1col25(0));
fa0st2col25: FA port map(st2col25(0),st2col25(1),st2col25(2),st1col25(1),st1col26(0));
fa0st2col26: FA port map(st2col26(0),st2col26(1),st2col26(2),st1col26(1),st1col27(0));
fa0st2col27: FA port map(st2col27(0),st2col27(1),st2col27(2),st1col27(1),st1col28(0));
fa0st2col28: FA port map(st2col28(0),st2col28(1),st2col28(2),st1col28(1),st1col29(0));
fa0st2col29: FA port map(st2col29(0),st2col29(1),st2col29(2),st1col29(1),st1col30(0));
fa0st2col30: FA port map(st2col30(0),st2col30(1),st2col30(2),st1col30(1),st1col31(0));
fa0st2col31: FA port map(st2col31(0),st2col31(1),st2col31(2),st1col31(1),st1col32(0));
fa0st2col32: FA port map(st2col32(0),st2col32(1),st2col32(2),st1col32(1),st1col33(0));
fa0st2col33: FA port map(st2col33(0),st2col33(1),st2col33(2),st1col33(1),st1col34(0));
fa0st2col34: FA port map(st2col34(0),st2col34(1),st2col34(2),st1col34(1),st1col35(0));
fa0st2col35: FA port map(st2col35(0),st2col35(1),st2col35(2),st1col35(1),st1col36(0));
fa0st2col36: FA port map(st2col36(0),st2col36(1),st2col36(2),st1col36(1),st1col37(0));
fa0st2col37: FA port map(st2col37(0),st2col37(1),st2col37(2),st1col37(1),st1col38(0));
fa0st2col38: FA port map(st2col38(0),st2col38(1),st2col38(2),st1col38(1),st1col39(0));
fa0st2col39: FA port map(st2col39(0),st2col39(1),st2col39(2),st1col39(1),st1col40(0));
fa0st2col40: FA port map(st2col40(0),st2col40(1),st2col40(2),st1col40(1),st1col41(0));
fa0st2col41: FA port map(st2col41(0),st2col41(1),st2col41(2),st1col41(1),st1col42(0));
fa0st2col42: FA port map(st2col42(0),st2col42(1),st2col42(2),st1col42(1),st1col43(0));
fa0st2col43: FA port map(st2col43(0),st2col43(1),st2col43(2),st1col43(1),st1col44(0));
fa0st2col44: FA port map(st2col44(0),st2col44(1),st2col44(2),st1col44(1),st1col45(0));
fa0st2col45: FA port map(st2col45(0),st2col45(1),st2col45(2),st1col45(1),st1col46(0));
fa0st2col46: FA port map(st2col46(0),st2col46(1),st2col46(2),st1col46(1),st1col47(0));
fa0st2col47: FA port map(st2col47(0),st2col47(1),st2col47(2),st1col47(1),st1col48(0));
fa0st2col48: FA port map(st2col48(0),st2col48(1),st2col48(2),st1col48(1),open);
st6col1(0) <= pprod(0) (0);
st6col2(0) <= pprod(0) (1);
st6col3(0) <= pprod(0) (2);
st6col4(0) <= pprod(0) (3);
st6col5(0) <= pprod(0) (4);
st6col6(0) <= pprod(0) (5);
st6col7(0) <= pprod(0) (6);
st6col8(0) <= pprod(0) (7);
st6col9(0) <= pprod(0) (8);
st6col10(0) <= pprod(0) (9);
st6col11(0) <= pprod(0) (10);
st6col12(0) <= pprod(0) (11);
st6col13(0) <= pprod(0) (12);
st6col14(0) <= pprod(0) (13);
st6col15(0) <= pprod(0) (14);
st6col16(0) <= pprod(0) (15);
st6col17(0) <= pprod(0) (16);
st6col18(0) <= pprod(0) (17);
st6col19(0) <= pprod(0) (18);
st6col20(0) <= pprod(0) (19);
st6col21(0) <= pprod(0) (20);
st6col22(0) <= pprod(0) (21);
st6col23(0) <= pprod(0) (22);
st6col24(0) <= pprod(0) (23);
st6col25(0) <= pprod(0) (24);
st6col1(1) <= S(0);
st6col26(0) <= S(0);
st6col27(0) <= S(0);
st6col28(0) <= not S(0);
st6col3(1) <= pprod(1) (0);
st6col4(1) <= pprod(1) (1);
st6col5(1) <= pprod(1) (2);
st6col6(1) <= pprod(1) (3);
st6col7(1) <= pprod(1) (4);
st6col8(1) <= pprod(1) (5);
st6col9(1) <= pprod(1) (6);
st6col10(1) <= pprod(1) (7);
st6col11(1) <= pprod(1) (8);
st6col12(1) <= pprod(1) (9);
st6col13(1) <= pprod(1) (10);
st6col14(1) <= pprod(1) (11);
st6col15(1) <= pprod(1) (12);
st6col16(1) <= pprod(1) (13);
st6col17(1) <= pprod(1) (14);
st6col18(1) <= pprod(1) (15);
st6col19(1) <= pprod(1) (16);
st6col20(1) <= pprod(1) (17);
st6col21(1) <= pprod(1) (18);
st6col22(1) <= pprod(1) (19);
st6col23(1) <= pprod(1) (20);
st6col24(1) <= pprod(1) (21);
st6col25(1) <= pprod(1) (22);
st6col26(1) <= pprod(1) (23);
st6col27(1) <= pprod(1) (24);
st6col3(2) <= S(1);
st6col28(1) <= not S(1);
st6col29(0) <= '1';
st6col5(2) <= pprod(2) (0);
st6col6(2) <= pprod(2) (1);
st6col7(2) <= pprod(2) (2);
st6col8(2) <= pprod(2) (3);
st6col9(2) <= pprod(2) (4);
st6col10(2) <= pprod(2) (5);
st6col11(2) <= pprod(2) (6);
st6col12(2) <= pprod(2) (7);
st6col13(2) <= pprod(2) (8);
st6col14(2) <= pprod(2) (9);
st6col15(2) <= pprod(2) (10);
st6col16(2) <= pprod(2) (11);
st6col17(2) <= pprod(2) (12);
st6col18(2) <= pprod(2) (13);
st6col19(2) <= pprod(2) (14);
st6col20(2) <= pprod(2) (15);
st6col21(2) <= pprod(2) (16);
st6col22(2) <= pprod(2) (17);
st6col23(2) <= pprod(2) (18);
st6col24(2) <= pprod(2) (19);
st6col25(2) <= pprod(2) (20);
st6col26(2) <= pprod(2) (21);
st6col27(2) <= pprod(2) (22);
st6col28(2) <= pprod(2) (23);
st6col29(1) <= pprod(2) (24);
st6col5(3) <= S(2);
st6col30(0) <= not S(2);
st6col31(0) <= '1';
st6col7(3) <= pprod(3) (0);
st6col8(3) <= pprod(3) (1);
st6col9(3) <= pprod(3) (2);
st6col10(3) <= pprod(3) (3);
st6col11(3) <= pprod(3) (4);
st6col12(3) <= pprod(3) (5);
st6col13(3) <= pprod(3) (6);
st6col14(3) <= pprod(3) (7);
st6col15(3) <= pprod(3) (8);
st6col16(3) <= pprod(3) (9);
st6col17(3) <= pprod(3) (10);
st6col18(3) <= pprod(3) (11);
st6col19(3) <= pprod(3) (12);
st6col20(3) <= pprod(3) (13);
st6col21(3) <= pprod(3) (14);
st6col22(3) <= pprod(3) (15);
st6col23(3) <= pprod(3) (16);
st6col24(3) <= pprod(3) (17);
st6col25(3) <= pprod(3) (18);
st6col26(3) <= pprod(3) (19);
st6col27(3) <= pprod(3) (20);
st6col28(3) <= pprod(3) (21);
st6col29(2) <= pprod(3) (22);
st6col30(1) <= pprod(3) (23);
st6col31(1) <= pprod(3) (24);
st6col7(4) <= S(3);
st6col32(0) <= not S(3);
st6col33(0) <= '1';
st6col9(4) <= pprod(4) (0);
st6col10(4) <= pprod(4) (1);
st6col11(4) <= pprod(4) (2);
st6col12(4) <= pprod(4) (3);
st6col13(4) <= pprod(4) (4);
st6col14(4) <= pprod(4) (5);
st6col15(4) <= pprod(4) (6);
st6col16(4) <= pprod(4) (7);
st6col17(4) <= pprod(4) (8);
st6col18(4) <= pprod(4) (9);
st6col19(4) <= pprod(4) (10);
st6col20(4) <= pprod(4) (11);
st6col21(4) <= pprod(4) (12);
st6col22(4) <= pprod(4) (13);
st6col23(4) <= pprod(4) (14);
st6col24(4) <= pprod(4) (15);
st6col25(4) <= pprod(4) (16);
st6col26(4) <= pprod(4) (17);
st6col27(4) <= pprod(4) (18);
st6col28(4) <= pprod(4) (19);
st6col29(3) <= pprod(4) (20);
st6col30(2) <= pprod(4) (21);
st6col31(2) <= pprod(4) (22);
st6col32(1) <= pprod(4) (23);
st6col33(1) <= pprod(4) (24);
st6col9(5) <= S(4);
st6col34(0) <= not S(4);
st6col35(0) <= '1';
st6col11(5) <= pprod(5) (0);
st6col12(5) <= pprod(5) (1);
st6col13(5) <= pprod(5) (2);
st6col14(5) <= pprod(5) (3);
st6col15(5) <= pprod(5) (4);
st6col16(5) <= pprod(5) (5);
st6col17(5) <= pprod(5) (6);
st6col18(5) <= pprod(5) (7);
st6col19(5) <= pprod(5) (8);
st6col20(5) <= pprod(5) (9);
st6col21(5) <= pprod(5) (10);
st6col22(5) <= pprod(5) (11);
st6col23(5) <= pprod(5) (12);
st6col24(5) <= pprod(5) (13);
st6col25(5) <= pprod(5) (14);
st6col26(5) <= pprod(5) (15);
st6col27(5) <= pprod(5) (16);
st6col28(5) <= pprod(5) (17);
st6col29(4) <= pprod(5) (18);
st6col30(3) <= pprod(5) (19);
st6col31(3) <= pprod(5) (20);
st6col32(2) <= pprod(5) (21);
st6col33(2) <= pprod(5) (22);
st6col34(1) <= pprod(5) (23);
st6col35(1) <= pprod(5) (24);
st6col11(6) <= S(5);
st6col36(0) <= not S(5);
st6col37(0) <= '1';
st6col13(6) <= pprod(6) (0);
st6col14(6) <= pprod(6) (1);
st6col15(6) <= pprod(6) (2);
st6col16(6) <= pprod(6) (3);
st6col17(6) <= pprod(6) (4);
st6col18(6) <= pprod(6) (5);
st6col19(6) <= pprod(6) (6);
st6col20(6) <= pprod(6) (7);
st6col21(6) <= pprod(6) (8);
st6col22(6) <= pprod(6) (9);
st6col23(6) <= pprod(6) (10);
st6col24(6) <= pprod(6) (11);
st6col25(6) <= pprod(6) (12);
st6col26(6) <= pprod(6) (13);
st6col27(6) <= pprod(6) (14);
st6col28(6) <= pprod(6) (15);
st6col29(5) <= pprod(6) (16);
st6col30(4) <= pprod(6) (17);
st6col31(4) <= pprod(6) (18);
st6col32(3) <= pprod(6) (19);
st6col33(3) <= pprod(6) (20);
st6col34(2) <= pprod(6) (21);
st6col35(2) <= pprod(6) (22);
st6col36(1) <= pprod(6) (23);
st6col37(1) <= pprod(6) (24);
st6col13(7) <= S(6);
st6col38(0) <= not S(6);
st6col39(0) <= '1';
st6col15(7) <= pprod(7) (0);
st6col16(7) <= pprod(7) (1);
st6col17(7) <= pprod(7) (2);
st6col18(7) <= pprod(7) (3);
st6col19(7) <= pprod(7) (4);
st6col20(7) <= pprod(7) (5);
st6col21(7) <= pprod(7) (6);
st6col22(7) <= pprod(7) (7);
st6col23(7) <= pprod(7) (8);
st6col24(7) <= pprod(7) (9);
st6col25(7) <= pprod(7) (10);
st6col26(7) <= pprod(7) (11);
st6col27(7) <= pprod(7) (12);
st6col28(7) <= pprod(7) (13);
st6col29(6) <= pprod(7) (14);
st6col30(5) <= pprod(7) (15);
st6col31(5) <= pprod(7) (16);
st6col32(4) <= pprod(7) (17);
st6col33(4) <= pprod(7) (18);
st6col34(3) <= pprod(7) (19);
st6col35(3) <= pprod(7) (20);
st6col36(2) <= pprod(7) (21);
st6col37(2) <= pprod(7) (22);
st6col38(1) <= pprod(7) (23);
st6col39(1) <= pprod(7) (24);
st6col15(8) <= S(7);
st6col40(0) <= not S(7);
st6col41(0) <= '1';
st6col17(8) <= pprod(8) (0);
st6col18(8) <= pprod(8) (1);
st6col19(8) <= pprod(8) (2);
st6col20(8) <= pprod(8) (3);
st6col21(8) <= pprod(8) (4);
st6col22(8) <= pprod(8) (5);
st6col23(8) <= pprod(8) (6);
st6col24(8) <= pprod(8) (7);
st6col25(8) <= pprod(8) (8);
st6col26(8) <= pprod(8) (9);
st6col27(8) <= pprod(8) (10);
st6col28(8) <= pprod(8) (11);
st6col29(7) <= pprod(8) (12);
st6col30(6) <= pprod(8) (13);
st6col31(6) <= pprod(8) (14);
st6col32(5) <= pprod(8) (15);
st6col33(5) <= pprod(8) (16);
st6col34(4) <= pprod(8) (17);
st6col35(4) <= pprod(8) (18);
st6col36(3) <= pprod(8) (19);
st6col37(3) <= pprod(8) (20);
st6col38(2) <= pprod(8) (21);
st6col39(2) <= pprod(8) (22);
st6col40(1) <= pprod(8) (23);
st6col41(1) <= pprod(8) (24);
st6col17(9) <= S(8);
st6col42(0) <= not S(8);
st6col43(0) <= '1';
st6col19(9) <= pprod(9) (0);
st6col20(9) <= pprod(9) (1);
st6col21(9) <= pprod(9) (2);
st6col22(9) <= pprod(9) (3);
st6col23(9) <= pprod(9) (4);
st6col24(9) <= pprod(9) (5);
st6col25(9) <= pprod(9) (6);
st6col26(9) <= pprod(9) (7);
st6col27(9) <= pprod(9) (8);
st6col28(9) <= pprod(9) (9);
st6col29(8) <= pprod(9) (10);
st6col30(7) <= pprod(9) (11);
st6col31(7) <= pprod(9) (12);
st6col32(6) <= pprod(9) (13);
st6col33(6) <= pprod(9) (14);
st6col34(5) <= pprod(9) (15);
st6col35(5) <= pprod(9) (16);
st6col36(4) <= pprod(9) (17);
st6col37(4) <= pprod(9) (18);
st6col38(3) <= pprod(9) (19);
st6col39(3) <= pprod(9) (20);
st6col40(2) <= pprod(9) (21);
st6col41(2) <= pprod(9) (22);
st6col42(1) <= pprod(9) (23);
st6col43(1) <= pprod(9) (24);
st6col19(10) <= S(9);
st6col44(0) <= not S(9);
st6col45(0) <= '1';
st6col21(10) <= pprod(10) (0);
st6col22(10) <= pprod(10) (1);
st6col23(10) <= pprod(10) (2);
st6col24(10) <= pprod(10) (3);
st6col25(10) <= pprod(10) (4);
st6col26(10) <= pprod(10) (5);
st6col27(10) <= pprod(10) (6);
st6col28(10) <= pprod(10) (7);
st6col29(9) <= pprod(10) (8);
st6col30(8) <= pprod(10) (9);
st6col31(8) <= pprod(10) (10);
st6col32(7) <= pprod(10) (11);
st6col33(7) <= pprod(10) (12);
st6col34(6) <= pprod(10) (13);
st6col35(6) <= pprod(10) (14);
st6col36(5) <= pprod(10) (15);
st6col37(5) <= pprod(10) (16);
st6col38(4) <= pprod(10) (17);
st6col39(4) <= pprod(10) (18);
st6col40(3) <= pprod(10) (19);
st6col41(3) <= pprod(10) (20);
st6col42(2) <= pprod(10) (21);
st6col43(2) <= pprod(10) (22);
st6col44(1) <= pprod(10) (23);
st6col45(1) <= pprod(10) (24);
st6col21(11) <= S(10);
st6col46(0) <= not S(10);
st6col47(0) <= '1';
st6col23(11) <= pprod(11) (0);
st6col24(11) <= pprod(11) (1);
st6col25(11) <= pprod(11) (2);
st6col26(11) <= pprod(11) (3);
st6col27(11) <= pprod(11) (4);
st6col28(11) <= pprod(11) (5);
st6col29(10) <= pprod(11) (6);
st6col30(9) <= pprod(11) (7);
st6col31(9) <= pprod(11) (8);
st6col32(8) <= pprod(11) (9);
st6col33(8) <= pprod(11) (10);
st6col34(7) <= pprod(11) (11);
st6col35(7) <= pprod(11) (12);
st6col36(6) <= pprod(11) (13);
st6col37(6) <= pprod(11) (14);
st6col38(5) <= pprod(11) (15);
st6col39(5) <= pprod(11) (16);
st6col40(4) <= pprod(11) (17);
st6col41(4) <= pprod(11) (18);
st6col42(3) <= pprod(11) (19);
st6col43(3) <= pprod(11) (20);
st6col44(2) <= pprod(11) (21);
st6col45(2) <= pprod(11) (22);
st6col46(1) <= pprod(11) (23);
st6col47(1) <= pprod(11) (24);
st6col23(12) <= S(11);
st6col48(0) <= not S(11);
st6col25(12) <= pprod(12) (0);
st6col26(12) <= pprod(12) (1);
st6col27(12) <= pprod(12) (2);
st6col28(12) <= pprod(12) (3);
st6col29(11) <= pprod(12) (4);
st6col30(10) <= pprod(12) (5);
st6col31(10) <= pprod(12) (6);
st6col32(9) <= pprod(12) (7);
st6col33(9) <= pprod(12) (8);
st6col34(8) <= pprod(12) (9);
st6col35(8) <= pprod(12) (10);
st6col36(7) <= pprod(12) (11);
st6col37(7) <= pprod(12) (12);
st6col38(6) <= pprod(12) (13);
st6col39(6) <= pprod(12) (14);
st6col40(5) <= pprod(12) (15);
st6col41(5) <= pprod(12) (16);
st6col42(4) <= pprod(12) (17);
st6col43(4) <= pprod(12) (18);
st6col44(3) <= pprod(12) (19);
st6col45(3) <= pprod(12) (20);
st6col46(2) <= pprod(12) (21);
st6col47(2) <= pprod(12) (22);
st6col48(1) <= pprod(12) (23);
res_a <= st1col48(0) & st1col47(0) & st1col46(0) & st1col45(0) & st1col44(0) & st1col43(0) & st1col42(0) & st1col41(0) & st1col40(0) & st1col39(0) & st1col38(0) & st1col37(0) & st1col36(0) & st1col35(0) & st1col34(0) & st1col33(0) & st1col32(0) & st1col31(0) & st1col30(0) & st1col29(0) & st1col28(0) & st1col27(0) & st1col26(0) & st1col25(0) & st1col24(0) & st1col23(0) & st1col22(0) & st1col21(0) & st1col20(0) & st1col19(0) & st1col18(0) & st1col17(0) & st1col16(0) & st1col15(0) & st1col14(0) & st1col13(0) & st1col12(0) & st1col11(0) & st1col10(0) & st1col9(0) & st1col8(0) & st1col7(0) & st1col6(0) & st1col5(0) & st1col4(0) & st1col3(0) & st1col2(0) & st1col1(0);
res_b <= st1col48(1) & st1col47(1) & st1col46(1) & st1col45(1) & st1col44(1) & st1col43(1) & st1col42(1) & st1col41(1) & st1col40(1) & st1col39(1) & st1col38(1) & st1col37(1) & st1col36(1) & st1col35(1) & st1col34(1) & st1col33(1) & st1col32(1) & st1col31(1) & st1col30(1) & st1col29(1) & st1col28(1) & st1col27(1) & st1col26(1) & st1col25(1) & st1col24(1) & st1col23(1) & st1col22(1) & st1col21(1) & st1col20(1) & st1col19(1) & st1col18(1) & st1col17(1) & st1col16(1) & st1col15(1) & st1col14(1) & st1col13(1) & st1col12(1) & st1col11(1) & st1col10(1) & st1col9(1) & st1col8(1) & st1col7(1) & st1col6(1) & st1col5(1) & st1col4(1) & st1col3(1) & '0' & st1col1(1);
-- END AUTOGEN COMPS

z <= std_logic_vector(unsigned(res_a) + unsigned(res_b));
end RTL;
